PK   �n'YQ��  �b    cirkitFile.json�]M��8��+���@�_`ݦg�}�iG�F���PP�֌,�J�v�:����*I	J �q\���U��|� �<m�ߪ�t��V�ߪ�n�Y�(�>��ŗ���j<zZ������m��i������x������f]��SS,�Ҫ�t�(ɲE4�t�LQҬ��"��j���q��t���e�ǲ�����Lvz.;��N/����N�;���#!�H�=����#!�H�?-䟖�{B�i!���Z�?-��O���������i�5QRfYd����Y��*Mk�7��A�;���<�V�b��o	Ӭ^䋚t�y%E�F�̪(�����zV'Srç�����O�/�6ږ�U����i�*����䝤'��������_OV&�)WdO���U\F�|�����,Q�1�-��ʩu������'y��dFEE���f:����EyU�Y�͋�,"K���2u��]i�J �~f�Jpei����բ��EDT�(�m;8ΣjVպ�5�9��No����|:]6�(�v-�x"��	�!p��������P��������z� �����6?��hQU��%x:���ף��&>T��4����p���4�K#�����+��^#��O�/ZX���)�)v/x��/��'͏��6?�D��O��%X���6?�様�޽�)���4?��G����ѽ����4?��G����Խ�9���4?��G��T�aO�{Ȱ2X��kѿ;V����be����W`��G�����_�{������P�"�S$p���M�Qu���8萢��0� V�����5 �@�	�"�ST|�O���� KAKncٻ"��C��(�F�``)��Z�8E�H�_)ף�`A����8E�H�_�أ�`Y����8E�H�_5ڣ�`q���8E�H�_�ۣ�`���B�8E�H�_Aݣ�`���r�8E�H�_��cy X1�`�H�"�S$p�갛@T�KW{D�O�>��=KH��a�OWK/{DC/IB�I,JB�J�Ql�O����(���)8E�����UkJ�)�S$p�NQ��o=�֔4XS�H�	���{{T�)i��$N��)8E�w���:XS�`MI�"�S$p�����Qu������8E�H��-��ȶ�iَ">�vG�����n�����Ҿ))p��㷦/�g�Ym�BO�џT�g4�� Q4$J��@���($J�b Q
�@�Ű�0�%	C`�0�0&�	Cb°XcX�Ac0���b�a�ưXcX�1,��,u�Di8\TJ�J���w¾4�ka���J�Di�K����?J����z���K�m��Z���K�}�m� ��~C=]\uK-��@���Y���W�7��{r�_�zy� ���%���	"i�v+ɝE�Q�H���!�Ǥy�^"L�?iãn���"�@�[&r�xT Ҡ��	<*�9�ܜ�4(i�X�
D�eZ-�1�G"J�{����nQ>�'�@�AIsxT �-���4(i��
D��E�
����[DS�=
<*��W��
D�47R�G"��Iஂ���r�7N*H+B7�c��K�a��0zY�"��
>,o�f6H�K�0ٌY���"�n��
�^�=�vֶl�ǂ������ǫ�7LBc�&��H�a*� y{\]@xÄ4f�����������7LNcV)��H�a�� y{�b@x��%�o>,o��6H�O�0i�ٯ��"�k���q��W��k̨�d����ǧ�w�
S���a���� �|X$�-k�>2 �Z��[�6Т�a���}* �|X$ް�i���q���טq>,o��6H���0}�Y���"��k���q���ט>,o��6H�/�0}�����"��k���q���ט�>,o��6H��0}�����y\gBlC��1��l�k��՜f�/��Ԝf]=��꼷=�i�Q4$J��@���($J�b Q
�@�Ű�0�%	C`�0�0&�	Cb°XcX�Ac0���b�a�ưXcX�1,��,6��G���`sy��6��G���`sy����ȣ��K�9�<
�/w�lN#�r����4�(��i<� �4訇� �Vn�i�QaI��[	`N��
D��ǜ�t�p0�AG"J�cN��
D��0�AG"J�cN��
D��`N��
D��ǜ�t˫���4(i�9:*��`N��
D��ǜ�t�80�AG"J�cN��
D�E?�Ӡ��%�1�AG"�"��i�Q�H����Ӡ�"��H�MZ�a��	L'$o�9o�T6�V6�X�S��ˆ��� �i�a�x�4�A����`���fܤ�7L9$o�9o�x�MZ�a�x���A����`��Ihܤ�7LE$o�9o���MZ�a�xô�A����`���iܤ�7LQ$o�9o���MZ�a�x�t�A����`��Ikܤ�7L]$o�9f�
L_�&-��%+0}m��}�4�a�7i��E�����gN��� m�i-IíIhQ�0�Z�>�9<,o��6H�>s�0}�����"��k���3����׸I<,o��6H�>s�0}�����"��k���3����׸I<,o��6H�>s�0}�����"��k���3����׸I<,o��6H�>s�S�oc������j��.������r[�O�r^-���t�]T��Ç������W��A]�a@)-�(~㾡� ��K��y�%Zn�@���!��Ixu]]�O�ϻ�'��
���`=D7IXM=d��p5�#n���J04$���������;���������yCxt����p������o��7���v���ڦWo�KoAT��B�
=!�����n>F�]�y' �y'�����s���Sy��3y��	9m��	7��}~^�_<�_~���!�3�~^.�v�S_���%�k�����Dx~*<?���7��)��2��$)IJB����4$)IJD�2QK���c���Z�D-e��2QK���L�R&�L�����x�.�d�p����b.�KX8҂p)�]��P}��<ȶ�h{V��.ؼ��s�.�ź�6����c4����n����W�Z�v����͛^�����E��wz?kkQ<��W=�a�02�;N�
���˘��ƚ8c��5.�!�T6��p����3�=#}�/�`�)*��t�:���AQ��Ǖ�"��u�:�킋AQ���q�"�#w�:�Â�AQ���M�"*�W��L�Ń�(N����A��Eݫ�����AP��q��Ń�h�L����6�Ae�I��2��;�=V�BP��ڽ�l�.Eq�3g\<��_�I<�E�!@ʳ�5b�D<p�+x�����L�\�A�<�+x$�:� �BPz�Y����X��2���އ�H��p�ʳT�h	�[	K��@�,}��R,:7�`	���Y�̐�X� n�� ���K�hB���%@g�31�b)�I|����,j8K�A�K� ��y�1X4!p�>�a��*čw�1�
 �8K���K�^�@�D�]W
-`�8K���Z��_�>S�b �j �r �z �H��
�(=Z$�&�R,���Y����XT!n����
�����J��B���%@g��b	P��}-0 K�*��g�+��
qkZ`@� U���zW�%@ⶳ��,�8K���K�*�-e�s&�ܚ.�4וs�`�9�F�o���&��¹[�E����Ç����:� sEu;��Ga�~��r��&�f�O�F���H�-���Z�kN�=�ȝ����Q㴤�ڝ��ڝ��ڝayt��o8m��'�5�=!d���	![ot�"�| j]�NS����ڇ�cz�zG���������f|��=��=�;�}�o�,�u.m�߿�W��uta5�7�
:�v�[f���.��|���s�ţ�o�tm[̷:p2��	��^��{�� ��Y�r�+���]�����vu������C����b~(9J���x(凲㡌ʏ�r~�~�8*�!:U�x9��t���[�r���h��7��r�wl��̾�Yn�K�8�QN�ҋ�6F����BOߕ�]5��U�ˋ�����ɽ �P3v[��{��b�ɤ8���bY��z���Z�K�k����S��/+7o��c�r�ܬm�� :���O�J&�1ũ��n�3�cJMUE]��&�>��8����Re�9¾��j�k.B㑝�����(d�2m�K�<tt�]��i��/��UuL�v?�'�E9Ʊ������]�5��M��@��v�c��7V륲&��x��țΘ�N�o[�"��B�f����T��v���3�9^��I�4���@�<�w��Oѝv���3U����6��t���!5)��DWN��ȕ����9�$��W�9$�v�G��2��vq/7�1^��.q�H�!�i�����0�vy/7���]�p�l����:����Q���A���؆p���5H]�e�2׉$������L���E�Oj�[��S;�^ǅ>�z�����^,7/�ۈ&�$�ϥ�Cma&q��L%'^Fj�{������/Fܤ�Cb�#��}"���,���Hj>SuRyG��j�R]�G��x=��z�����z�2z�g�vJ���3)��kj�Z��qh��vcWʊ\��l�efR����qK8{�$�}nƯU���1=]ဲ�Hf9��>����G� fm�5֙-�!�8Mhb��{�����4w�����X���:���0�L/�*)���j�0�1�a����*�Mq�����	�D��9�t���}d�4��c�n��^�t����Q\�Re���7�}ӧ2�����Y����颜/H$)���;��4c��@�z�l��i��rU�-w��r��u���쎎G���g������i�F�z^/�+��������O��ȣ�ڽۃ�j��r������m��}^n+[��}��X}.��u9�?o�?��ޅ�fg}y*��z��t�jd�s=�ϳ�}ʛ�gg��+q�v6+(�ha�Ѭ(�B�NY�"�C�\gv���!#kll�d��c�LH%���ԛvi�Ύ@�+�hl��;.��\0k�J�CY��&��~�D뢭�="���y�h��X�G%�![��amUՎQb�s�2�=h���B({�*k�9|����}8*�!��/�>�����+J9�T-~x����V���,�/����"7��q��{�GG"S�����h������/�?.�C�U�&X�^xB�E�&����3��6�����f�޿/����_?~�8r�������ͨ�s�}������qL��={쏮����|�lu�I������7��u��oG�,'/���]sH/5��P���^��v��%qL�C��X��H�>ߺ��`����⵿��y��wX�&���IQq9&�� �N�4eJ����7����|0��eJϧc����8��Ȕ��k�,Q=_b:tHOo���E�h�a.�W��Z��N�S��U����?���ś��U��q�H�>���X�� C<��Er�a��ڕQ���xǏ���a�(�3�(��N�.��v:�R�B��փ��Z��D`:�Ni���r�h!�IN��
�J�	Tز�J��?u�*p���mW�t����EԿz]��<`�*����(l��P���Jԡ�����s!�Ou�q��Z^u�;� �M�Z��^�;7�:̋t���L�n�I_�|���—s�z"�l�!'l��<�s���U y<��L���7�sլMŹ�;�6c3��)V�Რ	z%[�9��c�);��*rb���Y.��7{�^w�,U�4����g���f�/3����;�ˋ�E5�*��,���͙�sZ�vivZ�]�7���r����{����r�6�YV���W-�^������?��;���c��v��j��k��o�O�oۣo�PK   �n'Y��(��8  �8  /   images/12674a71-c981-4176-a988-13f1272e71c5.png�8!ǉPNG

   IHDR   d   �   ���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  8kIDATx���T����������tX�,�(HS�(c��5�ؒ�1&�3��&�F�1�?1Ѩ�1��i"(�.,�l�;���o�웶�]��|ٙw�}�s���<ߘ1cZ����&�x<��z���K\\�466JKK��=!!a��f���f�w||��{���!x�#��1��|>�< �\�r���>�v�q���͛eӦM2e����dܸq2l�0ٹs�����	��}�G�ĉ���J^y�)//��=�IIIr��'˜9s$%%E;�0ٺu��q��.�E�u�(<�]p�:,��g��:9##C$999�x�m۶Iqq���Yd��=z�̜9S���Z�߿����K����g��C9������'//���'�0s:T�-[�_�y��Jee�A<�~��f��ٳG.��2Y�~�����KlϧO�>2`� IKK3g�޽��555!�A��Ғ��w�O��Ө(P�6rݺu�t�Ґ���v��an�U�J�ٳ�lٲEv��%EEEf�u���Y����3�\\��� ���s�]�}�v�����3c�p�n�4i�2��Z���^�>r���J��/6���gAX��t�0ax�R�%J9�t�$(u���Pޚ�������_���:�\��B���w������a�\���ZxFvʆ��n6���q};Vw�%��W�^�JAAAȯ���S|���c�����#	z��!cǎ���z����iJ�=�!v�#F�xAW��M�� 7ʶ}�����o�'�|R=�P����
�%tvn1+Y������� �畕+W�"L�n�,�e���V�Q�������ؕ�;,11�E�[��r��p)�*�B	��-�N�����P�W���9~�m��N�ͼ�_�כ<���
-���?�8O���h��TU�.��w�q�lۺM�9��y�	RUY%wnO�
As��>عc��=�9����o��V`��+������J�,^ I	>y��G���e��r�7N�Q#�ˋ�?+�e%���$��		�fa(^���_���%�w����7r�5ט�7��>K�K6� H�6;D���}W^ye��gϖ;���S]q��΀Ҭʐ��������<�w���eM��*�q���Q�Ƀ�Յ���&3$>c��dű�;�H�lʢ��d᧋͹��\I���y���/iƙ��v�_�w�<5w����J��������7�IrS��Iz��́����n��{ｆ((ʶv*�W�=�c��y<�ET�3�^8X�A�W�ҴZ���:�h��47���5�����|��/���S��رn�(���o-N�#�:TD{P$��߷�rK���.�j�>S[[kvKT>j�js�bn��|<����5��Zb�(��s�D��Ǽb�]�yc�ӑyU����<+,�9cΫ�dT��?Z]ǹ�����;�4�n��V��+**233�#��i���|�8��$:�#���A %H��<T� ���Ȋ��KmE������"i�x%��@��;\�S�Ϯ�x�i�\�y� q���)��=���|�^�'i=�IF�A�OT6�����2���U��%ez��U��KL���C$C?]��MQ�G�EM��Ç������޽{�sss�a���)!��Y�Ǒ����=?p��G�e���u�1%T��Q5���]��SZ�S|2�~)���J�����LK���ee]��|��t7T
 �-�d�s7If�Qr�ٿG���mPB�{�ϲo���'�Jz��뽪*��I*<$���Ȁ����؅�����d�+wI��)2�?��l�����3Y������Œ���z�U5��a^�T��e��ߓ���"m[D��[�r�jY�R�}II�T�6��a]��t���O>	�!2����������<�4��q*�.S{dȼy��;J�/QJ������L헱��K��s�qSJFZ���`�������u�����oB�C]���RQ�.�L+�Aj���ŏ^#Ǐ��+�"#�$9)^�A�U�2��5r�_~*{t�#ξI�g�aW�W�H�����#��Z��m�+����3��"��d�jƏ�"%����ܵr��W�ލɘS�	��V����by���� /��1N�����0���s�ƍ1-��7L�q�5*;??�:%�uF�c�~���F�t�l�ʽ[d�?����)�~�̙�A��_��dמ*��'��8Z�N*W^��,zl�L��{%�N7kX�]@�ؚ�BY��������՗�nvqCc�46���3H#?�l�����e��"�}kP��Ƹ�V�;NO�d�+��;gȌ�#���IWs�ޯ�k�3S���'ɱS�ɅW>*k�H�Cg^e�+7��P9�}5V�}�,|d><�-�!!  
��+d͚5F�[�X�s�GV�p�\|Z/��w�HUu��`���x|�Kj�z��F����˟�8KN��aټ�e_g-��Y�>W�x��?#U���t����X��#�u�����o�>C�\����͑�+���#�}N�+e�[䞟-'��_��o��]R]� �����>SN��)5Mr�n�� W�����Ø
(F(EVku+FQ%2�V�u�r���l�XR*��U��g���푕,�Jk�fq��J�F��x����صߛ"���w�a���(ݱN�K>Tb|��Pb����݉�e��WL��zD���}^e�;�͑��r��ce��RIJ�Ib�W���o���
��/c
�ȅ����T&_pgTcֺoX�����m�H�ٴy�"����2u\OeK�RS�h��#E�o.uv���2E\��x�����c&��?,������
"�UVP��C9�l雗��v�Ab,ئ�n0��:i�yґ����[~��RY�M���z�{?}O������ҝ�7r#A�aR������Fe��N%��H��
�%�>?�(�����!��&+9';IW\�Aۿx_���K���{fF���U[H���2�G��f)��kŋA~Y�Ab4b;i�A ��/WeZ�N�8:b��F���)���Fz�<��&��Z�+��jw��8�i^��=UR_]*��i��ϙ ����M ��� i�	RV^�ȑ}5F{q�0��y؆�����o�x���vC�r�Ttb����j�So�[O�Yţ�L"R�qd�e���wX��7G�����;�c�9
�)��l�X��I��'����d�`w�d%Ii�#GXٰ��D'�V]S/{�5J^f�!�X���Ȗ�k���#���Ęf���� nϾ��̍�@�y�{J�^�r��CU��5;ο�@�����/��+�T�iI�Ĕ���q�All!�66�	՞�gw�1I>x�ߊ�:=��	#G6nq��p��~=�)�͖��G��[�ad�{�)QJ���I ��d�V�]�!���n�2/ZV������K/�dvq��18��6�\� �3D�y��ﭒг@R�bz�;
����	a�92HTb,̶vJ��Qr󏐵��ǞY&W\|LP�쑝���k8���T�?�}�����'�EU{q`�6N>xs������q�!�8v�@e��Ab����:o�ߒ�䌨;�Y-�AGΔyy@ޝ�Q��rQ[�<Σ�q!�3���(�W-��!3���"Db�˗/7n�~���D���G��)SU��N���~�%2lH��x�H��X}i��F+���*O@�Ϳ{M���i��g�Dod�^ϼ�N�_y��K%;;U���V�-I�NB�x#7�r۽o��M�2튋̼�1��<4���W����z�����a����Ӣ��IP���R��$�3j�s�q�ع�M��(";��w�5���1��s&ʇ�+T�M�|�=�6�䆟ɏ��K.��x饚;���o�+�z|���6K&�^�lV�k�1o�ae�)�����1�R~z�q�B���ei��?�#/,�Ȥ���80ٹ� kښ�"9���W�LQ��@������a���r������t�/��q0�]��u�WO��ɓMX�
�j����c�k�-�!~��������-?��L84K�A��(��={kdgY�d�<U�~�ʪ҃H3<<�^�g��e�A�O7���]��'d☞2����k���5����5����Hbz�Qm-X~�
�_���~ ;�����O�}p�Y�#�z�� o�U�e���s��e��s���B��!����6�*�.���a y���c.�����TVmZ!�%�ū�+}�9jȑ���� ݽ��i$e����Kzn~б螷��{����-�d�ƥ�֢�FcJ�/��3ɸ��m��H� �9Vr��s6�K�C����Stޕ�p�j�_W">�aه��)�����&\p���I��w�.��]Ch���hH��5o��o��0ZZu�f��p�sN�d�%�.��1��*蝘�Gz���~BH�ə72rɽ�:QrG��6GecD<�1gވ��y�b�~��!8q���®`G����x���!?D�TĘת�!;"rq�o�і� �yc�3os(��ɶ�����,Q�z<z=o������jYhP�����/���Ӎ�E�	~~��a)R�v���E����(q���^��� �|w`�d6R'h�[�*B�6�9������!>���3���o���  y֬Y&I�"DCT_~?��3C��_~�e�k|q-��{���>������<���Ki�A�cSe���ciA�x�bg��xꩧ��N$�p�Q��裏9�q�Fy�wė é�hb��8
C��;��c���ůApjR���7K�����p��/�ɲ���D;�7E�Q����^��J|j�7�oSF��!}����/�-/�چ��d�z%��(M���)��֔G8;էc=��c�H}S�|��"b��_r��Y�I	q��Ty|~��'5(�N>"KR������A���2���*�|��s{��Kf�7��U�9���	y\����Izr�؊Z���b|��+���D<u|�Y��,,1�fGI���N��u;k�9A�"�oR|����OvD�����+.�
�A���� ���Y�Z!ߜ��hۊ��Uef�����Se���^�j`�D�')�����^6�3��=vH�D��mv��\T/[����2@L�Щ���;����ʥN�N��}�y�N��t���Qį�V#��$^��6��������17��=L���k+�̱p��),k�:�����|y��r���ʱ�3ewY�4�[��D�����d����g�HB��7.5|�-Z-�,t2�T-���|;fJ��i�qf�r:�Z�1��}�RX��K@liu���b䎹%R]��w�V P ���c!pM��KG�׉���qeO�yڮ7d��-�+�T:�_���JaSd��dx^�<��^5�[�`��v��� �����)HX��u;k���c9A��� ����<�v,�\e��x���;K䝏ˍV��/'�9�^�Wf�a[EM�k_���%�D�n�wV���"�Kuek�(c�`��݂��sXЁ���,�3�$O�VR٨�ϰ"V��χ�~����nWM�N��0&S��y�҈�rK���ݶeo��M���f�F�o�,��Ň���O4i�6ށ7��؃0�X �6,-
�@�HeQ�Zv�a"��.�!�Peez$H�Z�ŕM��R)�j�0 ;��:/,n��}q�>٧c㾌;_u��=�g0ySii2x�`ٽk�,��m�)�ѠN5��gL�8o�*�^_Q�\H��=��A��פ��}a�HGE.���ms��	b�ymy�!x[c�X춋��Dbˬ}�D�����t��ҩ ??_vn�&K� �A�u��1��'�Hz�7��dm�]'��WF�q���c᰽c�
 E�,t�
b�]�z�!�������-Y�dI����s�1��t<QE���铝 /-��� PO�'G������w�����~wbY�<�B��p��4�����	��������5t�Eň#�����)�h4��?hA��x���Z�I���Q���F�N����ފ�#GP�H��[��t��T*�\x�&�Ǉ�E���_��C�Ô��q��E���)=Ϳ�T~���)Ƶ�9 �;i��4)S�m�����~���:*C��
� ���Ͱ+`Q�k�_z�%�e!�����,N��ɥ�^z�����T?��F����k+Je�jZ�(˸ٱ�Z� ���6��țE�dD�d�^�a,��D˲�������׾&�<�1;(4� �Un �$\�_ a�wךh��w�E슺�f��o6!QU��d�aCᮓ�6W��?�Q#���F�ފƮ���$�m�ԩ&Q���g�}V^{�5C�0�C�������8bH�	}���Mmz����V�I��ũI>��iʆ>X[a��l6Ao5 14�-J/��U[��;�m��� �J�޽{��ˍ>����4�>EV{�]���o\'9i�&"�Ya����A�a��_W;y��FTq°tc��7u���� {�Du����!�	'�`�`v�]�$p�� <���{�VY�&h�oeC�BeƤ�Fi@y���ii�.��B Mz �%�<�Z�*�P_A��A�����e��bΕ�P���������p0Z/o�ʛ[��<��kd���6Y9�,�E� w��/� 6 ��&���o��8Ot�kdA�,�Tm*sd��4)��aCh^�J5�c;'�Xe�ʭ5]j��b$U�Р��H
.{�A�zx��ϝ �bx^rH�Y�\�E��l��=tGʝ�4�U6D���I_௯,�)�g��66ICWʐ@�������3�qKM��?�|���,+V�~G�xx�	D��xB��q�/�P)o�Ժ�]��į�@Ö�u2�"��+��x;�z�+wrb�a���W\a�	���'��~��"�����J ka�s�8n���W��eJ�W��H�����yb?V�w��&��������#yJ�:��r�9Bl�8�!h�C�&|�nۮ��pH��SO=%4�a�!*A@.>({�UWy\�=�9�m1(��x+�A-�uҨ���+6ε�a/GI3�E8��8ix��O6A�-E��dO�!R4�C�����VXTѵZ��#���$^d	�N�������V�ߜ�D3f�0:5�0J�8�7��_C$W>/����T�;4Sm�����Ę�qy��p�z�if�%H�� d�'7���:�Ⱦ�f��ۘ�߻:/�P]�~�_�n|Ʊ.�&x��G���r�6Y`�jS����G�L�/5����$&����� KA��1z�"-Z�
G��;��T%J/բrt�3_a�"sW����~9�2�_����u4v����+��X�:;�o߾f�����i��v�te��5��v��`V�*\�XIZ�Wv�8�`&K��Dg<�jXRhB?4U�	�l��7���j��
l/i0�t蛪��jv��Bm���׿6��/���}�٦0�̰�o��4}��H9bB]���#z��o��b�X�P� b[F���S�e��Ϫ�C)D�<�'K�&��OV{�n�z��ޙ	����bR�
.uv��nM��I�g��|C��j�W���Թج���׿�e���v�i��B���QG%O?�t�	`���`U�$�b4͇��Ak�l��3X��d��&_������l�ߐr��#6E�Ly�G6=�N���~]�]�Kl�&�Yw��	P��!�C5��&b2ā�ݸ���y.���Ξ���,Аȟ��C,��!ҕ�Z�Y��C|n�CM��RGf��6� 	v�8���Ů�,rT[3Z���O����t�R�ԅ%�ǧB�v�DC 8qb����:a��r���,-�=�fţ1���0��`m�0��cL��d��GC(�� ��"�q���թ@�8G�?���r�uי������T/êº:�C��
���O7�%���af{���`2d @T�'�1dՃ�}��mU����O�el7ۢ�g��tY��p[���SM���|`ކ�]bm�zWc��b��`:��7�鮩�
���������m>.+�,D��hP�T��)kPA�J��v���#�EL�ú�dk�ݠ���[���v�,��+�m�(+((0JS�XY��ّ������{g���a'~Za�%���U[�=���j#kI�ț��V�1��p�WWB�l�r�{�����$�6�j����Im�u�=XS��E�z�hCMK�aSM��C��@�	lu׉���k��ӛ����x=��=jQ7 ��x:�[w�6_yp(Z1��	p4v�mj6�W�.��'O7V�b�I|q_"�'�����&>`,�i�B���iӦ���~!KȘ�-f����9�,�]���h���� ���y�xĿE˒�������w<넁8��w		t��w6��-�Ƹl�m-+���&����T�v,��]��] -�^cx��e����i4�g�ظ0��}&?����,�lMp�E�����F�W>�L�vZ��΅��.M�ˌ�n�y���Hqe��+�ND��c�>����}Yx<��ᮤP�`����m�56BC�dkjM]`�4L���� ;X�''���J\�<�JEVzs��ek�]���B���D7�K!$���3�L�O"�c��H�ƽ�lm'#q��d�*��,ͱ�!�7,����	�9pRw�pX<oر�.�}�!dH@&�w���z<�|�ȅwה�5Y�!������RS��a���\��0�.�<ei����.�/9o��K�/�$�{�P���4&x�ǂV:�!G�H{Ƣq��.!��{m�_�I!� i�x{�����n��p��`�I�t������ԟ�����$�ט�	�o��¿��`ߤ�m�����E�Ŝn$�PI�h�Ð���%)�qR�
PA(\�+�և8'�H0;���$�C�~xW!���2d.B��¶b�V !|�&E��>�������� ��XI�����C�����o����>:S�\P,q.����lA�Ӄ7��X�ZSx,�R�w�{�9I��V�Ww�#�����BXԨ�,z
v�$��w�$������]l�F1l��-D��LS�X�Dd�2'V���Ǫ�k��;k����'c��I<c�;������~�9D���5�6w��Pv &y衇̿�Xz4���<�yYT6��Wl�1�8�:t�|[92� C�ߴ�0v��Ϧ�'Ȋ���M.�g���Tn:�B��?&~ī��P/��îx����N�,`[!�݀��7��w)E����1�4P�+?2E`{q��V�k:9d�U�_[Q�dǻ�b��|-�f$�� �S�F>�Ġ����f��զdAc�˟e�� mX^��d�����.&��O����|o�Q�ρƌ-S���QwESk��n�#C'���Z2≭�0B�o� �$����k�4��x��w�I�c�G��`�;���R��-m��Ml�D��_�u���pv��:+�DY��
���"���h��:��v����������� ��u[�P��@nG�u%X�XW;�ŉ��x��fnl=_[t�=�6���l�. ��8a���Z�C�䴁g<�wSM���l#zsP΋��`�0L@*�M"�z��
2
Wms�O|����A�;���
r�P� �]���%���	V;�(^V�0L[�X���ɟ��'�$G˾�
����o6�YQ���j]�:����,蟓h�������^|e�-�}g��dD_��Ѝ�������JJ�z�}YV��\d�8��sx.��7��Ұ����~����\�gN�a�uV�W�\]n¸Ѻ_��N�|����f{M���;&��,V?�E����vc!���j7Q�=�����o�&y�^(AL��D�)�yn��R�~��=eцJY��ڴw�uB�W��Ū�� �WB㯊�%`��*~9���i��<�m�s��`S�_~�! �qd,��?��pm)V8ķ�e�9O����������:"K�_W�+��$���J0)A�+�X	QB�`�B�:*9���f�,��)��b�R����#�Mׇ�n�[��|�?��O�;��E(�`q������t�����R��g���cOd�����،Z���C6�ݽ��=TV-W[�*��}��D6;��d/Z-�*?�<0<� ����;T~yzaI���_Hn�(�nvRLA6V=����-���AHV<,���u��֭w5X_�o� ��c�1,ş��e�������'�:�EJY�J:��^��Vk�(M6�G��B�2��S"���� �2L���r8lZ~�.���~� �����w�qH>/� Ų6��|��̙3M�
q���7&?�	7�tSTyb�NrA/,�ՂgFXP�s��qJ����%��#�#�ߑT�����Gf�U�+�7Jr�	(I��%��v���!;�`�P�ЮP����?���L�ܝJ�*Lw���p iu�4bqr�DZ�-`y�[�a�õO8,���+��-��>IF��;�p'Ũ;hXoji0���x��z������`Kz����TиPy	\a�>�q(�/�����ch�A	 ��Z�D;��aD.q�ʭ����h0�!ׅ��?���^{�r���{┅�G40�l#�V�uCa����E@��� ��|�»#E4����
{��z�3�zDT�L���J2(�z���`;`��4�[*r��⻂�c���M��n��CU���8�Bk$����b^��:���z�T��[a� ��L�	�/:Б�� ��K%p��!+��HU�_��2 ��!q�����u�����!��C���i)��w�)�AI��\�3I�q�v���I�&9��h2W
�;݃�CwH�dAr=2��*$X��U`;ʡY��G�>��!������ �d~����"��[Kq���x:�Vo4)�MF�#�Q�I���=g��4+�a\���z
�J��(�tw�sw����fL�PB��G�駟JqQ���^'�a�+�Z��m����~6!��+`��+���o;;�]A(�gzp)���np�Y�29܆; �0)u#���P��kdO�Y��Y��*�b��7A��7�4�����r2����<]3cL���-�����o�����M2�n(sx�����3UgD�#A��X�$~�Z��H�:ݼ�1�0�L���	�$����.uH�)vH��5F���D9�= ٰ)� ���ļ�n1l� ��d3����߲i���47��Vt��c���pD҈�ҍU!Z�7Д̨�^'N�)*k0��`��w֔��v��N���v�!m�	�����闕�0Dj[��rt���;�=���pʑٲdcU�1\ t����-��&Y�&�3_W�+ٚ�E�(ma��6iҤ��B��
� =)@ H�0����n4��`Y�nք���&;�E�����O���Nt�O�"�.�	fB��K�`��IT2���w^0Sc���t��t��-�u��K�J�k�"�	E�g�u�>$<��Nkw֚RU��!Ć@Se�T ��^�:�N���;��|�ȁ4l�R����f�qh�x�E���1/z�V����ɼ4� �V���0�9�͜��e1���6x�(c75���cu��7E��B��9�F�H�!�$<P�jGյ��!���n���������=���Bڏ�3�˻���\[~C�u�RW�}Rp�p0;{�ؘ���i�iJ��h�!��.`�3�kk	��t������ç����������?Op�G�6�ڲ�X8�E;��S�ۉy��sQB;�� ��[�����ilj}��RR�Ȥy�����벮d����Om�\[��VbFgǒ�F��X��JQ��,"�L|�qm!x5�$�KCRRR�^�DO�T����'��r0��Ma���w�3�y��k�KQѮ�;����l3v��n�3����W_-Y�Y��ܹQ�Hj=�~�"��?�P��|�56+;K.��"s?�T�_�|��m������7�a�<l��n��D���Jq�[O����9��2���*[\ �b�)E�DxVO*ՁiJ�F�y[NN�T��Ew&�JZZ�uw-�7��ǻ�yw�;��n������ӷ��y�Y&��M����7jēE2$?_�y�9���/͑x �X[�y�̙m�Yބ��hԿoU�?���[%*�&8����Y`�w�!+����(׭7K,vɐz=�Dmm�|ec�&L��OG��A$�G�p��	�| cC�h�� ����x�� I��v|B|̱�L<)QbE��=

Z����>�r�s����}uʔ)�_}�U�k���)���AN�Ȉ�
�ڮ\�T}� ���Z�J<F�]x���|9!�r@q�/E~�4ü뮻�:]W�lYү_�Dr|6�DiP�<r��1 ��C�@S��J�B�)}��:P��ލ��ڇI7��~o��������L|^c�������<�a��(Q�Z�飼����u>��]��������q���j%H���>��?m�,��񇑛d���J�A,��:.-���uXEQm�@�䣧���i~Z����t��ȓ�L��4�o���L6M4��L=�p
�yْ%R��H��k(!�B zø���j��`���^�'e��z�=d-���%�j9<i.] �c��c��l��p��ז:p�v�9�����c��Y�<(7��"[�6\z��6oR�۲cG�Z�>b����a��ٺO��k
��L"GF�3��5k�.��8����}�ň7|���6x����{�rsH �M��U��'�b �?$d��(��\��O"{���N��'�"��߼�̂bAd�� D��o�86(�����bR�k3H���hK<0	h������f{�M����L����?_����h�����s衇>AT�7I�<�0D��曏�gK�(Rv��:CU����SSS_��� ��I�2o#��DA4��JҘ��~���7�
�A@������a�}�"�.�}B���� =B�O���l�~b�7�t��7��A�%��6���x.�3�-[��3f܊������.**���c��`^;��IЭ��^��:�c�٣ǲ�s����۷oϡg ڃ�E &q1�R�~�l��ްo�D�Õ�g�,�Y�f�����E�O�0��)�'�	�#��Bj/���XA^��:���[шY�j] ��g�x�\�E�\嘚�(q�����ڍ��T�w�����>~�a�����n�՝oP��	�:0U���"���^��ICYE��lKX�;c�>����<^[ K�=���3�!|�q���ܰ.x0Z	�x�qӥo�L�x�֭�`ڥ߻\�u~��{�9�d5����e�`��W]e
1�O�S2��P&M�l�s����:|�OԶI�{O5����ȸ�ɾ��ED���1c��{�>37����S����N,Q�fԇ��6���@�=	�S��֣U,l��`_��
?묳̃�7�Y՚�.�f��#��;��ew.fơM��Z4��-��m�b�y�7�P&Ƽ mlm��a_[�w��X����^����� G��>3�S�e=��S�>m!Da�^�ν�xFp�BR�'!�8»U��X�p�Lȃ�'uoyV%+���ʰ�`�Æh�ikYm�$n��p  �@2Id��؍n���Jq$���������ޛe��ܯ
�q����]�=Hp�柬~[�a�"c1��n$�k�FN� A6���^�wV��31��@�� '�m��9��]�| ��j��f���ժ�zN���w7����hv�U�16>p�B��&��}^o`�/0v�~�u���h8툽��� �u�嚶ȳoR�����[�B�t�uy�1ʧ����Tu��3Ϥ�؏^|�ŧ��8�t�6�f���c���o��\��+���cC
�u���=��L��e:�P�|��7����M��`��f$�8�U��� ���3�x���u�H��={v��D!�x��Ǔ ���ĩ����(!c�{T=�V��y%z���_�W�}г�}W�ࢋ.�")Ĺ�+ڃ&���UbD�E0G���� �`�灻/��_A��A�|E�n_���W�f�A�|E�n_����[�V�Ax    IEND�B`�PK   �n'Y8�w���  ��  /   images/54656ac2-7b78-4fd3-b315-813e86bdf352.pngt�eT]ݒ6�qww���=����7���N$xpw���!���s�����������%O�ڟ�eP	A ����*�A���#���'@��,��)F��A\R&�	ܥ��՜,ݽL\-@^^^,6�vnf&�,N�V'�� 9HNRL�;�軗7��@G��#WX���&$2RU=
�(�h�OLR���
	B�X�*�>�z�hP��2���H���;�G/��Ga�������0UD#�� �|y)_k%�E�	n!|�Q�xH��:o�'
�󊳡k���AV��Ehl�atܽ�V�}�-£�z��4*�����R��[C��sN,�4����t�P��P1�s��k�a��[��9Uӳ��$ceoZ���Hd��nD�N���z]`bX��;��n>��v���*/2��Ю+D�Ѕf2g��
ZU#��*�*�Ɏ�$�r\�gq+�R]�P��blz��r"�V�m�BO���N�J�Ӕ1>��Ptǟ��.�;���r84(#!*&S�����C�,�g�"��oá�l�mI�b��k�}�*[�:���rF�չ&�!O1ogX���@*�n��^i���KtW�U�,�p��d��v+�)tpʊ��мb�!�2�L��uh<�V?y�M P��<�	���?Sby�J������Hb��<խ:9�c��Qv|З�͉�c
�:���9�	�(���)HBOT�����p-��b��A�Aa���b��HȣqH�_�ۃ�#J��s�'��L�	B�r6���ul4{��x��i����=8�O�\QF	A�|�&�
>�9�Kv�mb�U��tbDev;ORq�`�o�Y����v�G�P��ˡ���h�3irq2��[�&�����l ��E�lP�骟Mߑ�J��2��E���b�RE��/��m�*�t�jz�Ƞ�*�M�'.a�+F0�6@��.g,S�P�xZ ^rߍ�!*���,�)e�q}	�z�"y�L�bTtE�Bs��$g.������u⾂)c���.ȉ@�F���t�>�b�XC��433�024rQ�I��ʑ��������H���L8�X�o\�8�qgt�w�t��|h7��*�� 	�O���bcP�����?y$S�>���Gb�gT2R��dܕ�u��|F�S`��Gz��)K�jY^��2��Fl������\���o\��8�\G�!�1&h�A�����m�"5��#��
�A��x���+n�<X~&Aڷ�cQ���V!'�졅��rx��}�Elv�4{↽) ����o+~i��K�#\�o�XF#��`�kL����0�TO-�;����"�Ck�������G�f����`b/ ��M��vgC�1|���Ou+�����ܕ�+nR�Q�1�.��7 f ��̫Č_��zE�E7�bc��v�ɑ�*�j	n�g�_&8s�S�J\Y`4`��J����g5%e����5�
D�6'9�eS!�G0���s��s�~�ԗd*@���%	� �[��J���0��)�nV���ݪ4UY$���G��6)���Tư�:�&�X?Ƌ�j����^�bs�7ߺ
J�M�i�S�ZV�:h�+zO�8�֕e�8DlF0�}G�SM.=4)r�1Mw�7��S2��Hb��)UG��>b#
��+0�B��6ϸ�������Y���Q�I��F�b�O��&�Y#
忶�&�A4Պ�@퉲��%�̇���5(b���(����7_�,�r��w[|�6�.$��W["3-��������'27DMbɥGg"yS�&�A(�3`qe�Qѩ�,?��ol
�Mb�KN�P�B��L�V���]Y �@�q"׬���p� �Lg�6gn�::$���/n�(��SʒĴ42��FE}VXD) QJ�|� �7�J&tQ��F>m�wzȥgg"��$�C�5	�:4iF��6/�$r��H{��3p�H�M���T���n^���ռ3 ��'C�h��GT�`�i��m�C
F7�;�V�~_f���BV�?�䪜B9����[�Ҝ������B�t���a܅�oV�ҷqi�t���a؅�%۬��/Z�-����:�B��/�֨�`q�{`9���@��"�k꿚��]�w�����C��0����$F��}�I����·�T��Qs�6M�C1��sX�n��V ��M��Bz�5���&�"\�/}Oto��#�ŋo�x4�3SHI��oWC=�/��@p�r�5�4�{f:�Yᖧ�d"�r4+���({I� | �B �!�{8��;�>��X�@;��Z,��l�qp�.����+����VR&���T�vL�Ц�ۅ���N�<��ٗOt^|g@������s�<�
�K�\�*���VT&�̿��,�F�ㆹ�-�P��4���:��Hy��e�=��f��Y���Vκ�f[j�!�Y<�&�}�R��u�r������V�v�Rݩ�����Ue�Yeu �d�R�{g`���y.�ddd��H��=�s����=q8���^�"l,��R���FJ�@?m��a\��-a*��T*ӛոe�:���:�
p�Z��A�f��T�]Hj�b���T@��1 �ah�i�d"�������3��h����_�|x���o��D�_�Ə��*>KR��뱖CJ�$2��v��fX�4�S}�Q:Q��:pEsR�#c\M�5�2k�̰�CK���������m|+'�dQ���^�(�r";E����;:���E�8j{�4Qsz $M�G�j�@�ä9�ˬ�Y	�׵�w��z�׾���>��h���;�Y'�(ݕ�Q�1gJ���,7f�O��g<C.��$d�� OǋG������Rl���f\m)ts�F��O���s��֥8=�҆�w6 ���]s�6���>�<|h�^��>�R�7.`(��a���gf\�����Rl"�V�D�J��Qh�1�<��֊̰Je��8��1�f��<�mUEH�'W�]er�X�A��hv���N��B9��vWC��i���N�12�X*�f�J���.�����ԩ+��N�cN+��KG#î�t���%��5T�����?�t�$CW�n	(��-�z�L�OѼ.��ƕ1�������(�Q^(}��v��I���(/�-c- 9�?y�]��ha?�R���+3����'�>ﰸ���d���z�a����^=�,�k� AP �W,��:O�7dcrP��8.^j�9>2lh�1�/	x����V
ퟛM�J�����.}񈌓�A"� �0Ɂ�^��U�3z���s������
�7���L������.CF���*�Ġ�Vc�儬vݔsZ��R$�2����`��3� g�)��� 敜�[�����^�3�<AL�J��r�ވG�G�>Ձ�ߴ���l)O�mJҷ,��v� >�z.Fe[$o�s<�F�,�xL��̾����}}��6�q	5����%��1��ŵ�4���=�HB��^%�m�������ԫ��~��ch5�՛�%��YCY펈��X���]�łM�&�"$�,��?�E��.����)��V���4R�\�nӱ�N���l��Nz�h77DȚ�����>9ѫ��߹���F��|�Q���ex!��z*�=
$��_� �y�tʹ�ǈ�Q�L	y�T�sNi�9��Ґ� �yM�7��)O;���)�̲�߽(&'�������W��;f�����=�`A�ivj�=KAͻ5����t���-P�G�:d�f`,��y��Wߞ�U l�x�;Eؗ��`c��(�q�ÕL������Cp5�7��q�E���4�e��F�R��P7�ݚ!U�h�Zz�c�����\���c��?v�cm|��������b^�_�zG��_���5泩�][5��q�J�.VVˣ��A��Q�~F���5��������+�,y/�N;�C1�XSLf/&�&�}��E���V��`��ow6wn��vj��ߚ̳ 8���[O���lԼ_F�%m�[y�U\��K/�u��FXAξ�S�^��xA��F��;��Ki�M�[U��۸#��j�$�mE=ul���Ҏjg�2hɶ�cA�%��eO���ǒg ��Ӂg�����U��մ�*�^U,�3g�{i��b�[����CvR3)��,��r{��i�S��'2�'�Q���R�>��j߻]��
���9((�=7�g�'�¾�V���BJ`^���#�J	-$Xy���	8S�wM��d�0��z�K��}�d+S��}xd�&��mH���@�0.�6�-ǭ��5�1G-,g@��s�boF��g��.����*D��+�A��P:�a�״f.��f���i0�!����J4�BM����JZ��)��?Ի� >f1ev���؜	R��؅l'=JD�6�lFnT��`�oщv#Y"#em�>���ə�*�
��UM_�_�2�pSC�Sx0��*68�]54_��� ��T�V����V���:�>���&L_�Ru��0�,�Ϩb����k�Բ�u�w-���X���Q���l�?T��S�bQ1#.�u�m���@�T����|�9��7v�ޣ2�P	���_X�/�R�j"�O��Q�����A�k�	)i�gR���]
�%?L�{��g���v�x����ZT�!5�%+��ɿ8�Z�~��"E�UW��$ ��+ʊ1�tw�X '�A�=�b�B�Uٌ���xl.a������|0	���	��G/S"kCax@��8�*�c���C|��	�z��7�7����� .�M����׽/w.�}�$���U�y)��>��US�PV�js��qe�dy��yo��<���L��F��E��|Yj<Z�b�z���0o*��O�Ƀ�4P;�v)�֒r��FTIw��y#�s2�6�N���"c��]ψy#ɟ���b���٢/"�l���۸����IS�0����a:?��B&)bl�M�<��pT?G=)Z���#����Ŷ��4ۍ�l;tXW~L�/7��볝�ϩ��t��_�"c; �������«�_~�_#�k��&+���>Be+�o�!mX�rX���x��hޔu)���2�B��H�ĭ�g�uë����j`��R�X+m��צ[�ւVǫ��:<�p���gtU_�(䋎��pP����}nMIj��?��L�A��n�?85�2�?�#��WQ1:��C&1�28j$�{tx�%&��\�8fvW�<�)$�S����:������?��S�h��#mx%�s���W��9�K�w�j���m�*�� J2R��vx!��!]���#敗�緵�Ƿ�����}W��o�!�#�x��/$�eX�-{H"�UܯAJh���<��hEq��;��OA~�]��0��ĢB'$9��j1��h}d��8���3���šg�:�c��W��[�A�$����}��]�����d��_?��"�o��O�y[�C�0�������Q���+�^ppMu`��7� hH��������������+����J�ץ!����M��'��H��S��?Kϐǻ���gI�1�kՋ���B�b�u�8�4R݈q����#HM75��Z���M7w��F�5���͌Q��^r��׫	�m�v�i���93�Ot���_��.��ٟ��.����8W��[�ǘ��(W�Df
��R�Ո�gL"C��v+�Iv���Ý�x"�{H;��l��9����R���`��ߩ�N��y|o^��ؓ�EҪ:�+�#��ɶ�
��*�K��Q;��8�1x��YU��B^¹���yR�a�BA��/o9��MqxW���>�@}:T	E��M��n�&��V:���g�_l�|0Q��m*�n�&���2���mSeR�&�cx�z����	���6�Tx�S��i��=���?������O
�bc��0�\8���L�"�ˋ�n3���t�O�,H�e�H@~W}͏��P��V�+�T`xr)�TOLb����T\���1 HWQ��ʃ}��ԫ�ŝx�1����y?|'x��.���٨�+�P���z1.�����>*L�,쯅�$~��"]O��N$���p��u����"NF5{�Q�m�O������MI����j�d>�u$9��|g� �h	�}����,-�\m���\ѦqV���M����/���7n'J)��Ts�w!�S�5��aE���\Yr��*�<�'O11�Pc&��ߜ�
K����Ǝ~��NB������Q�����@uf[߿�W.�`���Z�⤀�L$:����m��O���|o��{Ԣ�""8ȃi�M���á���wm������c����䚩��;�tr�e�Į��T�q���6I'� �4�u����2 W�rY rSin�����_9E0���4J���	v�'\5��N�ˠ�*�3(�� �Tߵq7F����B�'^-��3��������ej��RSv� ��>���o�M#1���|#.xmon��0=�3F��:�PE&��^BM~�������T7�&�fWr/9/�1�m������e�`YK� �.�k���0��]�+�#0a��V2�ZBh����#�cO��U���#!N�`¨�Tu������]Sܽ��K]Y��#�7�?N$��?����W�IT&Ҡ��63�j�yn)���$}�><熶u�ߚ���T��.���;7!U�
c90\��mx�.IM-�g��k1��w�v��7e�[��TL:�����!�+:��i3���8`�f��M&�VH 3�[�d��$}̯�"�, ��#w�ϔ�?�bcqo�)�QL�6�2��3���jԂ?�vk�i֦��ja�IM��qb������(�$P�N���Ŧ�J�w��M5�-p����?�Wd�C�o*����ȝ%��3�TjJ��f|5�m��,�T�w+X|x� W7���*�C����N.�8
T4��}�T��	����6�+yg����f�z��T�/���*F-zj��&sU��/��3I,/��)v!�|�ĺ�t�=�47�bj����k��4wv�H[9<�1�ރm/<�R`���T`S��c����b�3�����L��4�	5-��D��� �e�w+z=��	�N%!���N����j��%�r��O>N���8?�)��I,?3�d����K��j��J#�<4�b�h���L~��S
��\��v��
-/<=`4��i��7<l�*ڨ"R�,�r�UFU���n#Ü���k��;�D<��A�����j��} e\@��Ж�R�����Sh�lzU ��t�jv�ۓS&'�V���d.�	0��ߋ�o���}�H�c��ešA���i�U�����C?O'�ԑ�Lp������r+�P��5b3��g��zz���5~b���`���q���I9q�}
l��J0�L�r]E�1�c��᪓��?�=��o�OzU��s£�NG�v1\D"6E:���a�^X����D5hU��W��L��s�DV`�0�r��-p�g1�H{�@��]t���T�� 2U����5(gd@����K�*iL\}G�"����pQ�2l��+}&�Z���9lݠ���ʑD�|�Uҁ��[bed��Q��Y{ű<O �FU�:��	�?���c?��T��*�h�,I�@$7�'�eɪ�$�XL5H�����2	h�8��?n����o���Lf(�o��0�i�8�pK�^�����ȑ��sa$�B�;�?s�*A⃗�,����ݓV@څ[�(�!��wJ��|ğ����3���o�6Y�e��&���cp}��~�#����?ҵ�"�&�*��fETО}��tխ�Dq�Se!=��M2[ĉ�����k��]��y��64�Y뱱�p����������3��A��f&�\�$J�YOW_]��#��ʏ�t�)�s��3}�-��eHM�]�?�-��fkOn�M�J09���J�i9*���Y%�"��䵂ڙ�w��@wf�A|��x����j�H�rn�j[*�q�l���#jzS�B_��U���T,w��`�OM�ٻN��pC�C���	I:�*�,b���:Y� �C��<��PQV�=a��|'�<�B��.e�����a%�i��2w��]o���>�{�S��u�3�1�Nc���){��把g7�p���̑�	�B������Kc�����2�ʵ��v��[��'vz�#Ó���}8DÚ�k�z�1�ᰐ����Yko#nc��L���I���%�����h�v�B,5X���%���T:Ɗ���H�u�����p������!��r%H��c}�x`s�h|���ߓ��\*ɰ���Jl+��c�@
�|�z��f���-�&��]�i[L�!���`	���q�yrb��㘰�Q�C::����r���l*�!%geЧ5�f��O�=�;�mC�ެ����S_M�J2�����(�k�#�Ō���t�3�%��e�WG��
<�W��_U�s������c�k�.�)��'m���n`0��U���i`���/Nmp{?��g��no�t��\� Ǩ�F0����x�B8�O�B7;!&Nx3���1��
��>�U7�R�K�����R5��w��~>�%_��`�G���(z�m/-��pC@%��ij�H����$�E��OFH4Xj�J���A$���k~$�e�}&|3.�G��ʺ5?d_�{��z� �<����z$�\-�si)s�`v6_C�p���]^-8��h��yzv��{�[e��aq}���:�wvgW��m~�?l�do���ZN�]�ϝ/}�x�����ڵdM�m%�H:�7ܵq)h�MVk�>�{��t꽼�\"s.(%WLjU�j�֥VW�e@�K�9ޙ}��'�	f�|���-����͍���(�Z�s(�r�ӼA�D�����56v��9Ͻ�YMڈ�-@h��=�(K��$|!����]ܗ�ά����n&Ґ�`�I��~R��I3�ý�j�'^N��,��E���ƞ�I(����	"��� ??�����v8	-81�/�̎M�sj�,p�.���d���O��亜�D8f�����fM� O,�� �GAUϓ���4�2�0:���b�`�q��]O���]�Y��`� �E8�{��S��Yy5��l��e�)Q�I�։���3��+�b�{�����3��fx`lltY/�A���������zW�w~�Y=hn:��፛?�b~d<��:��S��u3U�m�U��G���������A��h�� +�~��*�F��4 ����J5'!������ta������yn�
e
�0��62�W?t�oQ.ѱV@Vn,?*+�c	�s��T)i	�����"P �{�-ݜ�c5e��F��{Z��mﻡ���
���ۀ L;L:O���}b���oa���{j�ߝ� ����dtB���eѼn7��pM�5�����{���Hd���l(��`�A��LBQMD�F|�iw���i��-�b]��͂��p��P�nY@���cT_�.Ywo�������jID�bh�y�Q((��}����h���}��� !Gۈ@�ȁV���C�p�0πɽմ��j��{�[�Ht�m4oJ lŘ�Ǽ�T�?�*^[de%y>ɐdS;&�'M�����t �W/ט~R�~�k��%�؛̓BDT�l{U�<�[��%�����i_ߩl
��B��E����zi8=kY�v��$�K���|ۙ#2���dɳ��i����@���;��� [L3À
��&��ۆt��5%�e����c�~ N<T�9y�Vo=+X��Ei���g#���\�d�9��Čp3�ݦp}e�3��>}Zy�N��z2f�m�c�~��aF�>KȌ��;�Κ�̘ؼ����c`H�ҙ8d��	������e����x�#�l�C`6�Ҟ���mWge���Z�CPu>ts���R�%��Ȧc��]�W��==��k��0X[=׮ߓ��N�|��+�^b ���o�Z_G)�3W��j�92�l{(詭��y:����n<���&{M��acpxHBE� �P*�&�����gO����q�%9D�Σ��
^:�1���,e?���LwCM][��iwD�v1<r53�$u>��BU�ҿ��_'�$\�R5�9�v5�7;}w;�m {���[���G{��nD��-���l�^6�:nj��ã��7�=��[�݈��ib�IERCٱJO�&�۩�.�4�-H&?��7RK�-����w�Ԓ�c�����(B��̯"��
�������Aۙ�0��먝���gdЊo�	�˪��U����z�·����c� �_\�k���c�-�2VpC��e
zo0�����1Ds����s^��Og:��f�h/�[��xU6���#���޼��ɞD�-'/H�\��a�l���}I� �G&�j�t�sK��g�bW��\#�=�� ei�΍��4���� Ʋ����VI(����u�f.	����I�����k}���ʅ��-�v�:��I�Ѯ����<����x�=�鰘#�����l���6�js���T�i�N"��W{��j�h��+�ox��̻ C���)ѓs�E�pzx�͝]��q��J��͙��{j�a���j��+��l"��΄.��+�[��9��s�*����P���]��z�s���fu�t��'�ZY�5��/4m>��$�.ӎ��`���{'�ǋY~V�R؛�(��O&}��g����N���ڐ/6�v=f��(9Tl�rXQ��� }B>�9�6b�sd@%��� B���y2W=�.^�^Þb&�^ԫ���Y��ؗ"�h�ܪf7�I����d��l֕��t���?�3��8S�����Y�󭆊��x�^pNJ����1��Yǂ���1�:s~�������@�����h�a�b��%�zh�a2��hOzfl���G�e��ӟ�e&�58��Z� R%v����-���$�O�_T��s�M�e�>�{���{��Q�7��h�9 �>..*✕=�[j&d�7bz\x��P��r$�Y������Ck�7ڌ��>uK��d��|�6�ǯ���������q��L����9Z����q�j[��6�.BZ6�_��\�� 0�콳6�������;�|�J������}y̞ޜ���ޟ����t
����Vj��'a�׈�BW����=�@|k9�4�W�G�,q��n��~ӺM@���~}v�EY�΁@�U����B��ŭ�AY��―��=�Ps}��V�m�E�3�����H@�����S~~˄�4��|u�խ��-�����Q7�L�fTE\�|9������� �*˻N�@�)��
�|�+˔��x���P�M���\��������6Na;���ĵ@$b���d��q�7n}��1�^���cBW�y�=�_�^絶����*���q������� ��ǣ�]x�� �҉��Z�>kN����2V��%z��d�t�󅹌���Y�ـd��<؍//�Z���A���v;�>-fUy���yz+��ܾo��sK3*���/�&Z<6�S4:�s�U�V;�����<�J(&MF�'_��n�&׋�ʭ@��?i6�������nk 2�֤�b3�>��
\P�\�=~������>�DG;X���O{E>_ �
�UV��@j�m�A�����p7-�������GY�q��^
���?�n/�\Q��Y���ڒ���|i�"C����/� k�C�6" 
���9�N򕡕	�8��IZ�x�iO��G��0gD���
@ț��޷@����^h����B�o���v����S&����!h�]�" �4i ,[ϐ�����{Y�qc�&[BA�2X��8�x{�!<H�'�zά�G
 4�;�r����� 5ҷϘ�4��j<y$�ueB�w��P�ԍ�p!&���ߓ�<Jb��^��R�ޏ'l��P��h�-'-�)�8]M �L4���ͬ
��?u�b+��q���o�̑-nAy�K#5S�a,�ˁD���鱃7Y��[�=��Lޯ��ָ��h���L����ۑ&q�}�[݄ɞ�Qvv<T��n^��&JF|�r����H�����Wr�;�h|��"}EH"r&�0H4�L~\����
��.�E,��v�_<��9�B�Q�8����J_~%�P�n�h��l��e�����gN�,ը�
�����.��w�����5&s~��P�P1{�7^�D�v�����P)����C$�������:R�6z5$<��!�~$�����h���[S��y���Upm�JI\��k�6�f��A�Ɵ���vF<�?��;�q7L�]�M�1��b�R������ŝk��V3���WR/旘��Ɍ`�jQ��J:�t�$A��[�8�=��<����Dc�z4:���O�P���t�/�>�.�ߜJ�ޕ�:��1�d
�i�a�,�����3�7�8jH{�,��.��=�v�GY�-{�ޏ���~n��5��ΠMN �4��z1=o���m�ZG�.�l�An�[������`�!v��� t�0P޶y������{|;n�
v�E~#�����-���4��[�?IO\�X��t��S�����\p��oHa�t5�b-Էd�u��U�:"�4�>�t0'�Glǭp����<���r-�چ�p4}�<a!��a�|yFu|��K��N��z�  ��n����>:Z�ĥ���b�M9����BL�\�������#�~ �i]���]8�ݏ�:r{��y�eN`f3{#ާ+���k!����U&�Lа}Z·:�5?Q0HqÞ#ޗ�o!�]FU��8�5��w�TqKq_}�	c	I�|R�D��&��_�l৕/���Om��w;d��0�wfKb�����y�(�(u��\��u���Fa�������L�A�\�_��jP�bPihX����k�!��I�y�eA�9�f[j�3%�_����M�T?u�>��ru���c}/:Bz��Q��υ3��=�4�d�g��0&��?�>m���FȌ2[b���6��6`���(����^8��#���l������۬��&__d�s��_��ӎ�٘*���oI��8M��,����i$�5#�#�� �c��,��|A����2Oӟ�&�'�6��,s���z�����/;�G���.�Y-d�}VHYݍ�Pg�Id+q�Q
�}���3��J2��F:弜�z;�yVU��������.g>�u���@�;r���L����,�ɣ�DԏM�Z;��F��J�IXb���cS��ɍ7�*�RX������+�X��Y�_��a����������|xg��q�7�u�c�~C�eY����C
�]@҄7��p�5�4���]}��lɑ��
yv�\GG?��fz~��*�Ts��x�
���u�]�k�W��Fч�	�Q�������W��׷h+��M�hftK�3<���S����7��|!��~�y����bIc� �v�w��cb�����S�J������Q�������X�Сň��XI��퇇$�߼H���~� P(u��q�������T�L����9�dm�ë|fUr:Q�QX+d�^d$���B����QX)�q�G�+rrr�J��x��u/�}[��!iD���[���KQmt"�Xͣ|��5��]���~�^nc�u��l��c0J�o<�C�����E�k~	�o0嚱{E�>�L�Dp*:j0��_LE>�Fq�o�S��fKگV��ގ��yk����銀޷d,' ���!�
m�37�^�4�1��8;��]rfd�:̌X2�bo	u�H����E�C ����&�2�2�W�uE�J]��\i)I�av�|=#�Z���ݬF���1��Vxh8��{�l������ޘ���������p�����f��_�l�� ���znl���A��C�2&�V���7+��!����f���9\��M{����-����>D�"��[=Ku�@5�i�H���7�8L����:�۶0���/.��3:���fޓ�T�D��b�e��[���~\��S����%@�����͔!"����G%����$z�)bw&�v��'ۆ��7�i	�M�T���"����c��jD������LF�F��
�!�4�[t���͐�wFd�o�T6��s���~���f�Q�I�s�����M�
L	i�G�Gٿ�T��'��ʴ��~r��ƟLw\�)����\uN�@���G���M�s���	�̥�M������[M	]\Y��U��d�2�a��$qv�� �<ǁݑ��
hV�o��(H#^X�@T�d��kl��ZW\G���\�D���Q�>6
Ѣe|ǈ�R|Ȃiߓ�_�Y]>�h/��I.��ՙ>�p�g%�-�5 ����g_���&Uӿ�4�(�zs�A؄���ɉ�Vpj�E1���x3�p%1����鈯��vBʅ��F&U(\w��|6a��IhDI|��[�1Z��D��i��q��}]��ߝ,�T�y���ݾy�*�7�*��n�F@�������<���ε�*�22��$~��T��h�s�&]E�Vo(������{}��
��o_H��.O�] k����DhF?�n�YRq8�(vn����0?����`��ƅ�"o�̥��cx���E�Z]���l����@.dd�)M�c���D�L�k/�\�>"Qa��K?6|��q����ff�i�y��XC���Ijq���>�Sg~��hr����ř�N�f٫	ܛ�ݲ��~�1�#��p$�yؾȵ�s�����d5q�=�,���t���iyN��Nj��tL�/�ﶵ���ɉ�e'�����vn�,�·�_Y��s|���~���t���{n0�c�����ŢR:����݂w<L��*�i��\��t~'�>Y��f�aPꔴ^*Uk!��|4�����@�v��A?G
h �����ͣ51���/x�3�I��h�_����7�*V+t��]����F�v�:OLM�}e�$�����Fv.�͒�O�R�<���u�F��㖩��?���h�6.��"���vkR��5�JYhh�5E�W�6Z^���[��)�	�_~���3CB=��9�(5���������� ]<g���������v��8U˕�Ӵ��{�nӺ��o}���
�o5��a���� 2�]�E���5P��cl�n���S�6_!V�}�#��bi�j�h��Vԋ�Qo��8�0㓲��._n���7��aD����C��1���ɱfM7n��k��;].j�k���#2 4q��7ȃ�̝2gM���%�G}3o�C&³j���b����I�Jb�MkZ�i ~ g�>e(�����������ҙ�7/C�Yd�~Z(5�7Ii醆D�*�A����]��X%9�E�Q���w�[�q�WST�A%+�-��/t�b��I��������^�8��X���L�{���EX����`�>�1Y��$���? 8�M��gP�����{�#���"/h���NYn����7�W�$hu�z�KN�B��N��� Ѐ��,l���f�b����gkV��5ӟ4���O�pG��ø��s#�����>����.w|��Q�LBR7:���O�Mݽ)]o������k���s"�ΰ|1:��f2O^�����H4u�zGN_���p�����Z�^�?�x�b��������v��`�<�h]$�89��o����sf�
��2|�S�zE�����e$/p���`��g	�s�0R�ĳ�{q��Ӡ���,NA�����ޯ֓e.uǹ��*����{���_K���qG	�2���eT#��|��Q��N� �3��C�Ņ����[S���hi*��8��L�
e��R���T����sV��3����j�$m�`g�Veۺ��v�R?�<����C[�5x%���`ۊ�pq���"ph����in�/'�t����{0>�����AZ�V���L� d+�4eO��lԨ#��^"��܏�ZK�7�G4�����.5x�Ά5��b}ꁋE��`ShQgͨ���-j�&��v�`VC�+���J��z��9���"�� h��F��Ӷ��D)亢�3�q�$<݀�5D�x!"w
>��+�.�H;�h��/�����{oCۺ-U�縯�q]XX��Rk ����k�ފ�������D �`���.�x����m�%��x	��>�["���y�ǲ��LW*�I4���I��!��)f�� ��G�m@ze	��(ح)��tX��n�cNy��Ǎ4]�?��sH��E �#V��t�Jr��z�/b	b��c�B��;��w���$s=�~s��*U��Sc�����!i�5�����2�;���^.ߏP�Nz�yE��ゞ��=[�9$��y+�y>}7,�mw@^ͼg�����~{����������>xT�ݺ��#15��1�߃K$cv�"�q��O���zn�~�������v�/b}�3H{��]�N%�{5�}������4'ec�L�H+�8�����!u*���)��_�NM6[`!-c�FW_ 
>wH�n>��Xƴ�j��3A&<��CI�G����7 
��D�+:��~�p� �=���,���={��[����0�%N�|���Jj�O< �I�\'V<r��(�p�z���&~��S�e��N���*�xo�*�ǉ�wg5� {�ۏ�'�|�d�.�sc�q�Ƿl�����j���EAT�D���R�w��+H�5� *ED@A@z�%�BT��tBh��Jh���A�s�c�W�=��R�^k�������=�,��jG�Sen��S �ۻ,�K��3�N��|N�!|,�|$�ΜcB�褎wI�7�i�$E/(	��q���������U/����l��mM�˕i���r�)�H!����]ߡ,�-R�P�{�{��{��k�ec�d�4:���Z�~��?����G� �0�Re���d�
߬�SE�#��G��L�X�W��3y��Nڒ^�P&؞y��/D�L]W��ȣn�>H֦���aF񎩯/qB�	h�:�?K���U�O�g���.�nkH�����³�;*�2�3��a�!��G�`8e�5�)�-��q�������u#
��I��`�y�:����t�)Q!��S��N���k�5Ғ=Y]%>r�F����=�q�\��l��h Z����% ��@�I�]���!����	��"���!�6�@ڵ��@w���7�_�C:�M�&��-KFPf�1��!�n� =�A�ۋ�ҋ��Wyy��ӛ�p����5��I��8 ����!�D�����[Op������\���S��P��@���k_zE��I�n~�1]��lI*L~� ���R������BZ�x���p��>v�&�����ʒ���R��K��-�~�D�b�� '�<9��?��E��:'�o�����}��H�N�C�>}{J�F�iL��9��  p�Z�G���^m�J6�ӏ�e����؊�zb�4_�2������G*�.s�����}��0إ@�$��;����*ʎ<&d�g����[Q �lK��'^b�Wb�h�n0]�<�����e4���O{�:�^���I�J��5X�M@�GV��}��G��c����Z�����ѝ�N��BZ����B�	�|�R(q+z+��F+}ނ�M�jaQ�d��U�|^��g?���6��z��Y���מ�M��<�� 1h[��xu����e`����)BH�$��٘F�r1n���)/�=�qu%XC�+^2߭�R��v3K�1Cu>�=��J;Mͻ��Q����ܹ=��)Q�\�!v���SE�ξ#�gs����R�T�k��}-�i�3_�n7��)T��B�2���=N�뒼���Pza]v�m��ۛx%������/�o_�Rpd��X�ʞs{��@B��ok���N�:�J�}����Cx&�|��5J�qN�) 4�P�W�����[@��(�>WD(jd��.�)t$���Y��T��3�)%|��b������
�>MFq�=U�>~wŤ���1�\AZ(B���_�O
��x����ܰ�i�WPT��n�s�ܴ��#n�Q����!�n��۩xܔ�%�gT��Ǘ��s���H-ҫ�Tgʲ>.O����Q�a���VC=x�{�T�5�jc\��ٍ��X�-
��-[N�6x�ΕbeHvs����A��8-���	e�k����f	����\cD���P�*�:�=.fT�޺k!m�
�F��-l}�W��~��	���Y��#[�ߏ<b���ŉ/	�Emmԛ��&���ў��eԨ|��)�r�_�A��b�a�-RSkH(�	�GB�cas1�A;���U~�0���utr?�\^lK'�`C��wi�\�&���{�dAc��*S?�9����f�w��,J����^>:��,l!�8yC��<w=������))3zњ��:�l�s��:0��ycm��cB�5|����<���7k���b�ל؂�.RK}�?}�]V�����kr�����9��}���d�TT0\��x5�k�g��c2I�ӽۋKK��gU?������\Ն������*�Ŏ^��r$�zq
7vt�UyoF#�RR�wM����I����{��A�C���h��a�J�[��":e�����=8���T���?8��2%���������'r�ˋf�BZ3��BZY�h}�|
��&8�>S�.�o�ͻ���O��'������m}5�c�;X3���m�zb��9J��2R��o�����|% d�xq���_^��y������{��^�'ĿxBxI�⛇2���H�L/>���#y�����jh�~���%�z�i��$�j+�'�פi��c����N�io2j��yCM�y�)&A��|�U���U�~RH�cF�����=$U��A�����$	�����!�ǏWu5�_D�{��F��Ab�8�t����1�1�]�������s�2N����J&�B����'��4-e�*~~�וh4dF�k8SV�֖.oe��~$���v$T��O�/�R��뵠��gМ�:t�JE�Kŏ�c=�&E��i�LaZJJ�������~~Mj�"Y�)Bʱk#%�D$�?+���PX	"I���O��L���&��&�˙6V���1�k���_RR������������G?����=9�cb���ϰ�������y`���ڴL�~�q���}��Xf\mԸ�Sk�����  ���`z積1�=i��^��,,}�Si\�OĬ%RhR�t0�������w$���6J��PEͧ����'����V������X�ii���҇z�'��nP\����*�����3�����Cf�����9�S����k�����;݂�P-���4��O�'8R���Ƿtgc��ua~s�zo�^�ώ���djr%���au�gm�O�jZx`�^�˼����^��n�TD%Eȱp����g��(ی	+/���܄�h�m}��<�J�K����0�d�{L^vo��|؃�6d6�F��ϣ�����N=��ᾒ�;�F�$'����*�ǹ�a�G�5*
� �&�^i�Y���;9�>����4� �t������U	�G���/J��P���b�?��΍'�^�lPT���xM'{�?�ka����%�{.S�'[E��Z��ۛ�cy+L��ʵ�2��y�Q��ڇI�ݶzm���B��Q�Mo�X��՞�Rl����%竤b��;����0�%���	���;�̝�Ȗ~�e&���/���L|�^h'��ш�q�y�3|�1�  iX�z��\; L1 �e�̩ķ���71��qx��C&��_�,��wML����'���k?��ܨ�zb��J�C�p�C�|��#��>�8o�l�d��P�YF��wMsҞ=��h4!є�bY��棯�^X2�'m���a��dK�n�NJկO��t��ĝ�QKL��t���+��#�����"�7��\�L��%�� ��J=d��	�޽�@����Dp��14��B�>����_"�DMnWҋ�*���@���k��N&#�ʈ[�ѿxp>]��f2�)���DY}e�3��2)zQ��x"Ϟ����&@>խ^*�]L�TPX�ſ���~�w��łR�Wo���'�v�%�=�)b�׬ H���8����Q��j�"�;
�a]���nP\bb�EL��:WȲ\6Xy�f�T�"c���{�/
���������g�=b-YZ��ؓUX.��>��T��U:!��x�f9���DHL��6��)����Ʈ�:"����F.%jp�IG�d��R�&����a\z%�~e�u-�!����)�7�Xa�JGW$����e�P��&�FGǎ^��,+�R*$��Fo� �~�	f��J���<~�M�vd{E�իW�7���Ĝ�솬w���D\�1$T�	�L?~��)J�F{�1~��O�Z+T��j&�@yR��ro�G��臥�J�d
�j�ڗ��L�NTք���0 |�Z��H>���=P�"-����\*�U�k����;����N*6�P]d��ؙ�c�Qd�`�9;� �[�Q�֐u��S��O;%N�5�B�+[��Qʤ�� ��}\�yU�����s����Z�ms���cx���"g��3
O��t8'����@x���
y5��v��g2��Z��s�A�+z=��`�6�Jۮ(������I~��%H����>�/u(��Ih��ܴ)���>E���r��7�f�7�M4��3D4%�����5���)錬�L��?*���u-��q�"/�oF�v�<ο���\���Ԩ{8�E�����)&��*K;�����@�l�)���_�6��܌p?���.�H��0�}o_�'�������Pɋ�����j}$,ژ��_����n���G.Zݽ�&�s^X�ouР��855U9jy~=�F�yV�b��z��տ���zl�a����1k�[��k�ɩq\��U��߼�R�9?��df%�����5��uf�իWB�➞�x���#<k8���8e%%=�0����p4Z�:�B{�5?l���$'�[�&j��;��!i?��^���H$M��p	����A*T�â҈Q�mT�z|��GpW��L%����N�y'��͚'Tu���oJo��)�=:�C���Lׇ���M���,>4����~!����٨r@�@����|��}��?3=r�����/�����dYe�|�ʓ��C�O��	��������Ǡ����6�vj��㗷�5�{��Ւ؋�I-#L2A�ɡyMPr�gFщ��Pr���ʶ�ӂ�d��������?�N�!W��""��x�O �^&���|�v�J<�u�l�r��F9C��#����g|�M�۵�#�:��M����/���|d�����LÌ�|o�krW�w���z��>�:\����Nx;�TV�8�@<~�,�y|o?v�GF��������U����'�ċ]�Q���>3� 3���7�@�o��̟���D��Eb��ŕ7g��>D���@@P��X����E��`�V����ʛ6������63����C�7�cf@C�jt2՝#p��X ��x7ٳ~c7��1��W?��r16ˆ���3o�?�m�ZKL��*�����U��{ITm1b+����k���]|���Sp�� ��~�9�ؾ\�׌g0�������;�%����	g�UE��f�X��7��}�k`8��z%��ǧ�����r�rm���ݹ�oy��/�V+8�G�F}-7�0��~�;� ߯�V|a��4�+�z����X��M�'�c d|��[8�M�/��2�� Zெ���RN���Cq�!�/�<=Q4���.d�qOqv��+�>�_���>��R>�D~�$���1�GE,h��MP�����O��wl1���Z�3�i�� � f������V����y�?z�Z�U��\h��т�r�f7e�������u���q�[�5���O	W^^��a-�X�V�A*?�^q$.&F�3n�Vl-����d���#Q6�N��1�he�g�7�ǅQO�q���NЀ8��Y�;���69�n��z�ZQ>���!́G:^/���5�J�~nz��H|f3�mw޴��dSP|zc���KZ��m/����V����C��Z��A�b@@3	e���7"NɎ�J�˅��5�:�f_��߹Ɲ��5�w|��Jf�bW'Y�9ب�'�εz'����PΏ�z�d��74YM�*�:�܋�GG��"��+��mx2{��P�\̤�&H�4�"KS=�Ye�;�CIE6��ƴ���ҵ(D��C��H��JM+�e��:��+xݦX��9OL����"-f��@gBO?P�$����o0��"���������u���-)��wPi�ym�OТ���E%�Oa�p`A8>��	A�	~��7��P(�N�W�A�z�71�=��`6X�w2�f�BO��*	���Ϩֻ���]y#%.� ���VH�g��>,�|,V�uU� �[���P�_�eL�_��Cv^�h>�&z+��C#o)&�\[:o�3�6յ[XR����7:�5�=�ES��'�?[��`�Y���ܻ/����������g6 �52zL���^[��i�SW _�ݞ�O<���32?�8�p�&��D�&�щ�|j�scrv{@������QL���y�@Cu��G����ϿJ�/���o�)o�Y����>r����d���9�1�>�v��� j�����'�1�I��B3��Z;�?��@���m\�>����~J���%S1$���H3O���Z���#r�j��5*
��� w����V�.@�m����HVO����s�'�x��y{���=^r��Gj�U�G�"��}��Vv_I
�B��T�iv�����V�kQ��l�?E��i�[��QM0"�����1��̬�{3ѧ�\OaI�dl�$J�0��k���'B�a�' 4��))�)���]�X�)��w�߲��ON�|�@��?��Ly8C$IM�T�c1x|�3 �K5Q/[��N�����{��<v�%�uq�]]�o�܀���++�q�~$\~#!)����cO���홠�m)ҧҝWؿf�"B��6k��P��րχ�1��Wi͟�o]����-� ^ׂ=HT�2���^Ȗ�U������˼��ݰ�-.|l�=/�(59z�oJ���pY�ބ��������o]�(ص'3��ֺ����}�IB�RJ�Ѣ���52`zhH�TL�H��~�A�d��4�+t��+ی	XմT���B���[��\���cn�+u��mqwW��R���.��M�zg��4� �E��'�����l��Mtm~P�G�+����v���L��=�a}[����	SN���c�/��#�ӊ�y9����[-^�'�B�c�rNVc����xM[��%��!���.�7��3S���ӥtr	�����&#��=>VK\%���T����ƞ�w���W핖�E���P`�zHUȗ��!qK�C�(f7�Х߮+���9�a{?�B.��Т�@ѐ����U�2����uv*n�T���gJ��)��,�Σ�3,׸�2��;�ds�V�_>����`J�������w�7�j�e���>,�z�����+���N��4�(�z��I]f�S ������r�ʽ	쉶�i��]�i�댲�����rϙo�=�m�e�&#h���|�|�$�B}u&K�� ��٧B�뽖��'9u���ڕ#��s��r���]ɓ�����>"j�NQQS���Ŗ'K�V澷���tI�kv|�(>C������%$'��Sꞡ����J󐇛�z�N�	Ʊ�<K�ڼs����3N�'v������ַ����^�Y i�����H�`�����G�b�k:�:��}����\�"@�]�z�iM1�mH4��3�!��,k�Ԉ����b�_ִ��+�<7?�XCtޤ�ω0�5.��l"x�F��C�C���Lm�X̢���2w�8���i��^��>֬a6z-b�R8��d�gZ��Z��z���Q�jH��5���v8镳2ښj��֋RR�M����ץ��J�yp¶�{֮�^�b �.���7 ���O=�t����D��F��5b0G�$���y|�ܠ.-��U}����Y�[¨G��Y�bHz��K��f?M5�Y\��K��f'�������j�q p��C��H��v��K��j�6�Q��C�f��qP��Sm�d,�.�:ʘXs�F ���;�ؒ��ҽt��L�����)�M���6[��h�ëۿ���,\��c_��l.<�?�N�<��̃Tb�1�ǒ����ɂ�q1/���J䱇��tͻ�{�>c��Xr�X$˝ӌo7/on	�7[�� ߫����x��8�@��ZѷOƸ'�l7��`vR��G�P�5@f@��2�D�'6��X0�m�"O���R=Ǿe��R>:i�5�|\�r�%C���LY���y����m�-S[�V^e�*s-���_�j�f�Dآ8{B�˶���T��ĪϷZZO��k����]��M��*��� �wl��nc����5�JO������$����6�(�M+z�҂V�";���Ϡ��W�p/�d�?/�R
��ʿ��^�pH��+��*���5zd6K�	��iRe8�$l�Y�pD�O��"p#�|��CA����#T��1�C�)V��(1��Z7�upߙe��Ρ
Ł��1�o�shP����p�Gkmkjzm�z�����6��V�������5��:�3��j0���G!�1�����Ă����>�����V��������BN���K�C9�F�CS��j'�YD�����=U��z�*�o��f���.�[B�9L�~�#7�#���:�ܽu��Sr)���go���w���h�v�V�)xsʿfr�P���u�#O��v��5(��G�4~[ЪK�҄�T��xu�E�wWM��|6�R fs��)"�E�c�֏���_�Y[/�4&�|)ryef�޴��L�=d�`��A��=X�b�M6�W'>�n�>j64���P��@}�L��&��!�%t���
�}�����_C�Nq��q]G�T�G���{f��l	�b"��jc�Z籟�R'6��&|���>)*�zJ=��p/Ȩ�7���fKve���L�"�r������<.�Z{��ؑ�IR���A���>l��������6�% �r'����6�F�Lw�gm��<8=SQT�ez��\���QY���u/�Y�>;^��\Y��<�Vd^������4��*@�<u�4�[��	��U�1Z�pĺ��b�N)2uXF�]3e��Hm��=(��V/�f�n-ߔ��������n��6��:�r:����]ss�ޯ�o\m�'"OM{{�U��#����~!���t��%#�>�&�涘 �"��%�ٞ�������IZW�o@�_���XԹ�x� �1	�׹�ܼ��!���N; �*��A�>�j�B�<�9zۦ����+ut�>ɘ
۽o�-��q�����*�Dŷ�b��@+��)��K��y�[�/GQ׈WRS���x#�Ej��Z��㏻�����r��]Ex"#�"*�S�N�-�Ddk��g�#j�Ï��P���s���\�-���˴'ּ��tЇk/0���6�U��eA��>�s���?�9*�ϡ���;rh�.jz�{n���,�#�|��l�c5	A�o�
������67���e������7�p�	Uz�2;��I���,Y�=\WO�YEc�ײ�ȥ�C'4��X(��f��k�dT�E)��:r�i�nX�V��^�s�Q�����Hl=q�wz=Qk�t�
�z�P>�EA���:+�U��a�о�}��ﰠ���-�@$�����\��<9��%�$�s
��+���P��,�R�ʝ2\��0�}�J�f��Ipꨣ7��x�@�؉Y�������g�o߰��ի�S��hV��Y��=bZ�{�i�t�&F�K�/�u���t�3&��\b����V���W�fN8z�$C������#~͓�\��

O�~���<E/]	DY��P�<���d8i�H�|E���m��-A6唦Ӻz�^w��y0.��@�~��5h�`�@���VՍ��/�/6R博�����y׋x��#�3 ��͌���Vz�����#�}���4;�!c�R�TD)�.����	��-aL�g�^= "�y[��I	�Ҝy(+�z����d�Cl{Ֆ�F(�/_�7;r4M���$$��3h���1��L<u˧(t�oe@��a���ٝ��MZ�F��A�
ݗ�{�R�W�X}Ƙg�j��R�u��k�1M�A�ޯ�0_?Øz!1c�V�"���v)��?z0������oЀ?l00���'R�mҔ5H[���*`�~��>lv4G�1q�7L�叙(v����3_�o���u|��?~t,ț}C_, �sG핻��g\,ʎ��s�ؗ�8��p�r��&o��2/�u��'���o�q�T:zY��f�_��c���kN�V(��ijT�5��'�"4 Q��*���\�l�B�y6�^��#EV�H¯j�����g�Y՞���U��;����\��<�����]'q����yĩ����݌gsq�(�`�J���qM�MI,�h�N�ؗnD�Y�ln^��(�i�����PBXX݃\���b9����I��ӫ|$׶K&�3�\ba����#e*��7Vk*-5m2 +��}����fc>����U*f`6Y�"����)��6�Z
툅ו��/T0�0��>G:	z7h08%�Զ�)?�r���{�S	j��LM� 4?HW���`_h�s��I@��Qs���i1sk�Y�Y&\��}���2 ��(�pRDl�܋�d��r@6E�)���7!d����r�S#x<N��.ܽJ����0٨���j�-8]mt�(�Th�Nbn������~���}vP��-����%�Y�%]�� ��tg#�ܥ�-���Q	.բi��>߫���Z�h�d� vW�y"nrʱ��g��x�ku���X��a��%��Ӄ���%�ЁXTV ƇP�U�Z���3��h��얃�����f5��	_�E�V�t2�P{�^�v)��X�?ȷ=�r
뫷[,@ Y�; �T���޴Gդ%��Ѐ�;qУ Z�+ܓ}4J6vP.;9LAS#.S%��[����ljA�j�y��q]D�)�k]U�������79����|`���J:��}n�r��.ט��[L��CĆc�Fu�;�+f���"��aX�^�� �+��̩ʻ�'�� �g�8�4f�y˶�t�?�c�|�.i��(r�
��d6Y�܂�]��S)!���[d��M����p�ʖN=K7�Y
�8W+�n��%yLz��:�ϝ�����I�(��Z�$= ��k����m�q����X�1��r��ͨ����,���q�?��ȓǜ	Ks�|� Y����8��\Ir���U��J�3$�YЬ��$����('^����o�(�K�I]����x9��-��-&�e�J��[�������J�))���Z�0�+P�}��.��f@-���Gg��"�^HdVk��Y�|X�f��$k� �i;�Mk��OGj �9��ǋ Ӌ�%|i�\�UW$�?Yt����aZ�>�4p̕x�f�asҜ+��|t|)M�[B�q���o�|�Sļ��T/2�j�\}*���`RO/J�f%1���͛@��;�8����*����Ý=��wg�u�s1����f��Aɢ�n���.�IO����@����e�i3�e�ZX�����,,����%�cҦ�<��Hhn�In�d9�6`�z#�؂%�'È�-�F�7��ʫ/:��@��q�)�8/Ib�-(��:�J��_�o����K�#�!�uJ/��A`��vvIj��S���%�+Uc~Evj��d��c��ꌵ��>�t��2�����`����<Q0����`j�{|l�����zba]�E��!�:=�νSdKy�o�/:,�Ald 9�돦ٸnG��;k�� ��l���P���t��$����y!r�KƐb�yi�5���ю"��	a0�p8�u�ԡ���p���T�0��#�'��
��<K1=9��/<MJ��/\��^ �����OYn��o�����"v���[����Y���ef�\�u�}�l�A12�i�.-�t�g#B,ފ�pOdn%�ؓ�"u?������k��a�1���B�*�+���ð���
au�Y��|��w�5Tu��T]f�}�Jº�- ��N��L���/Tz�њk�^���O�{�%e���p�S)BH;% �<ۭ`5�B�S ����Q������mx�^ǉ�����E�3���F5�*�C}r����bC"�Zs'lȁq�LC/['��?+�u�0���Xn�:?�u���զ�Y�S\N'���e�2�Yv���F��n><^}���O3�Z��]��	���+'}�G�5��{p3>�Z�&{g�Z���|���mJ��^/�p;5!�
%�}�g�`�"�7��HgkÃ�D��Zk=��Zh}��OO�˫NL|T�뿙���������8y��+��.����k����u��AK�ˮw���B�3�t�y&�����8n����ϛ�U�&�����ǢN:��%xN	�n�%Í �1VӬ\�� Q_9������U�O�m_NGӏ�[�vB��mJ�^��@Ң�K�X�1����!��O�B�S���"P4��Z�O�Vf��R��{���*����ߢф�
�==���F��&j��;7X���#3�S���UK����gS��%yf��$CѦ�7����������\ � �W����ޙ�������A���c��T��z���_�vK��]ݐ���:��n����Y�(���k����sJ�rͲ�����t��j*MJ\\��[����׸�^�.|��
��6xic�����p�#kp����][�V�H|�^��]qau��R�-��nUWO�P5o�#o�zm�.P���Y�Թgz�Ɏ�j�_a�Z1��׽����u@v�@��������H��ck��W.~;K+Y�/�l��3]jg�=�S$2�D�:��+�I'[����H��S1@�ѱ�k#�y���7A� �@kbN�6��:���ϫI�F(��{K�q�ڵ��)vI�6>�<�%�?�'=�cz��܌�p 1�<c����l�K����L�Abꑁc�'[w
��5q�D�)�E(U��像�[3p��|b&�~'�r�GQ�g�{O_4��ċ��f��P䰿IS��W��ȱ{M�Cʟ~D3K�0�)ּ{ȍ��,:�'���g�Y�rzR��ԇ�6┍8�A���z���:����mJ�&����Zʺ�B~۪���=L:<*I�z "0�"g���oO�~-ɥfw�csQ3�DhOʰ>��KGX�`��P���ZY��m>re�lÏgD4�7,����0oee�Z޹Mw�2�q�,N#4���6�3+�����O;���1(���)��~v�C�UL�Cj��gN>�ݾ��}w��)y^���QD��L��s����D�z��	�������rS|m�flC��_9�B]�+��Y���&���+r��&8��ϫ�}q�q��Ag��a��3�⛱Z(S�����r��p�9e�|M`�@;`�?����B�Dg�w.�A2�d�,'�J	�e�D*��wbT*45��z�`�C�{ WSRЉ1k�b�#��zN֨j�g�R�ȮR� X��=5�ed�;� �n�?:����=x+�AU�h���ˤ?���a6��7�*���!o�lv0�ۧ
0�)V{�xn����%���?�.xbtӛ� 
%.}sAN��k�!������p^^���Į��EYC���j���R�7Z<?��:���QK#3��-c���}Ѐ�rM%6ȑk�� 7M�����0HR�`(�[�"�#���-�Ε%5������YU�K<��n���,ֳ�|zp�\X�����6��jOj��R_�/$X� ����eA�D'//<���$��l�#��ݳ����C��A�C#D�������?�qD[�A�����xK��k��1�O�է�̲��Ջ�}އQ�e.Q:�HJ�Lx�|`������oT%{��C˴>����%���6�Ꞇ<eY/μK@����o�&ce������X��i�,	m��k��}^�h1s�K�n�>��М�I�]k>_�$���y��&Zp�;��#�v�o�+�����p��0�`�=B����������qH]RK]��_>O@]��Y�֦M�ȱEN�r<qi�:��Z i Q6��lX�%`;np(j�3�M�����/ii% ����il�Z��b9��8�f=�4hD�����<���:����Ma���!a��W��(�л��gV&NEs�ΏZg���Ż�|�˃�шj<�:�U��1I�aH�퟿,���Ԏ���"��N��w�?���\�h�y`��Lf#��m�*�Q�^��ngq8K4/��������t���;���
��X>Q��h��JZ@&�y@ܯ������ӆ@�H\\���%'6���5'������)�D$1����!�v����=�IH�D�h���҃����B��q�B;rQR�H��=c��EƤDdo�Hz�.Q����\�A��N�[{�¯i�۞�;��(���E��f}��vL�^� �0$���!�z$ �O!�Օʫ�T�,
�Y
C^��wۀ���O� ^�e�e��b��/���m���l�l��μQ�L�e��Ņ�ZS�ev��Zq=���nR���x���ݭ}�,����� '�R���CUPb�ã�X��5�ئ7���]�ρ��m#=0s���`�������������s) �o�K 2��}P���� &i:�����j�p��(�媆m��m�^���̃�O�b(OB!�3�qV�] ��.*�� :����G|n	����h�I{ɻkn(��5�mr��i�v�����W`��,��cR�>*�k�'G�ڀ{��w1�r�kʟB3�s=��*w����� d���������
�t�y;mh����d]��ٸ��������-Q�M�Q1WH	�A�x����;�#E,�eDD��5��z��rVX�������B��ܛ'�'����w��V���}*�:io#֕���Z�A&���c�LV������}������.;�/С��K�}�Tr�8�.��7��M�L��(����'�vC|��#}T%�J��9a��H�%��{忥Z�Ԉ�Ă���c��ּ�[����	�`�Õ��rb`�^�4m5���&:�^���������7?�76�%G�[�m���i\h����X/0�E�Ը��D���y̩�ܻ�J�3:�2#�> ��Y���Z���j;DW����7�q��-��N�'c]x 8
��a:X !�(K�{̀,U�K9|ZI�$��O���8)��"��0�o��po~���c>$���E�H�����-p��^w���~{A�#N����ö���󢉭&&q/�����<�Q��u����C6���*HM�:��T��]Zx�<�h>���1F��`)��T�ڋ�Y�o�^|�u�I��<��ܰ�D^d�@>����c!�ί����r���Y:��cʒ��{�˔�=D��X�������T�[}�R=�" ^���bV�Y��~Xm����RD�0G��O���ަ�9�� �i��ვ�@׉S�n<���N������҄���/�U�ИD�NiȌ�}d�Ɋ_|,��1UL��@tF;'.��_��涴��8(Vz֭׊8u�<ꨅ�댙�Xq<n��Z�[0�XX؜�c��<8��V�c���w�*�R�@���2���~" _�
l8 ���_�%h�c �Hu��K����LL��
x��L��9�>?G]�xϒ��^X�X�B��W[<yF��	��*���I�����pߡW��Q��i�@���#�h��3��~�8�����P�jP���1ſg���Ʀ�򫝾%V�G���$�-��sӬOM7�p�q�����jL��>��AY
��?��z��"H����(on��#�|'���c	3��bL|�4ڬ>?�5S�eQ4��UTT�A��~��l��w]�z��'��mʈ]#��!~p�L�a�,��+�س��kޒ����V&�ꟀGiL�*�{拈�a�?���F�l�c�2��敟J����[��>:<�iR�&�P��e����4���99����&�0��}����������t�º�����T�Uʆ�MK�${u�Ø��@`�1�{J��U�&Z��٧�-�V�.ϳ��~���A����LNJ���M�M�X�1W�V�x�����k�Ap�có"u~��u��@7�M�,������j� }������s���=�Ԣ�28�#f� ��������J�9x�@�ğ��P�[���\�3i��hqr�2��wx���l~l�*KV�{���c/��,��F_�4�\�ތ.0�,��U����8%��I6�^��U��>�|�G��r����S�l�N�x���Fh��|�1p�*��X^�s�Q񊕈�=����	����\b!c[�����{���XU��2��v[�65�Y,����z|M�у��������`��p]���p�=�\!v�7��<"�C��}�<��ܐ�v�X�:���s��;���4�33�z�Չ�_�B�����=8<�1�}����6@���Y��x� �D-K��3����ދ���˵��Q����"`������ƣ�!��LK�C���{"O�m�҇���j��	x]�~wI�F���O�|�wן]�|!����+v����$ro��5��/���]
yCr{`���Y�I��9�˳��W^����0���|��2�o9�	�����D�B���T���7��iK_�t#�Kt��1{n�-E�O�Au9h���,W7/y��'�/=�����;�֋fB��u�,Ά�v�8��0Jy�T��ޅx|������'�q���r�IM����������*��t����}C	��I�H��[�~?���3њ��Q�Y�'�<��� �v�:go��W+��V�¸�<[JyZϥ���_Y�H�m�|fq9�b�0]�9Cȗ@�rUk��wi��U��SPý�����'�蛥=�;�B�		��x(��}	)�W���u��]�F��Y�k4���V|fu�}|5�ה�y3�sk�B������ ����0>���Ծ�v"a�󷫼��.-����f�]�u�C�����?�tS�
_����[�Y/G&�Yq����cPa�TA2�Ǫ�����ڕ��?�|���jT���.p�0弛5�P���q�9�[o�N̟��(Έ����~����=��3^���ꭙ�.�АKb"�T���a��w�����Ņ%;�\�LYB��"L�i��L潧Z�o�2o��8��|�*�ǁ�����n{d��&����}VV"����*�"j���+�����>�$XZV��s�?�96>��ߗ�2Um��]�:�,�%����������z�����c�/"*����+�:��(�� ���w柽�����y�tu��%��������v�����
�X���tp�[�'����7������n��:�PO���}+������x����Ľ�2��>�ۖ�ou!c�v�����{�!|�������M6�q�������Tj�Ԥg�Gm�������j�އ������CBZB��������K����n�z������l�>g�Z�z�}�g7Hg.��ұi�ӐHd���م}���=c�ՋE~�),ȫ]�-�W�u�NN��u��"8�h
��y}@���G�������X����IXO��JSF \�8�o��Jr,���O����0��U(�@��y��^s�T.�s�n��/S1�Svھ,gsqÛ�y{6��� ;�r���������c������X3�9��s��'�p�1p����36:��9:�F~n�jd���*�qWo&��nWp��]��S�+3��L��	�=|��]�>�-��M��]o�~Y�U�\2��)G����"��`���d��=�`oc����+Wc��O`|�<o��U'�!�� ��c}a��\�(��,3�g+h=���ɨ�L�I�w���(�k2�A��(b�FEj"�&T݌����c���F�ᱣ�cC��+K��4#�� b0nK#65���Ǝ����z���Ȟ�0����o^5獽C#,�¶�bP?	�j�R6����Ց�s�ҟ��4ᒐ�D��CJ*Xo�k����%�<$��Ƹ��+��(O�s�j6$�U�F>��.A�\s{�7%��yy�(�)l�=�B�=���=���y{�e-AxrG0�Q�����k�*��a^�]��f{��砗�ܪ~H_j�l����lg%7��oʠN�����]��~�zywhs�*F7�:��wh�����d� �ϥp���Dk�5w�I���N��N��N`�\�n/�,�-V�P��6�42���&���o;�	�GY��t;�y8#K�8�	�a���.��&ێ�_��<�ir�׊]��;��\!3��z�l���ptG��)rI��֢A
�
~g��VBn�B�F:�L?�/93�$;�����dN���@ܿ'G�5��7c�=Mln��g�Gw��Ǽ�����M^����S���ɴ$�+i<.x�C��u{��:p6� BC]��LBFBY���pa����y{ȅԿM�]5����[Ն�M�������4�#g���X�U�fg-ߞjܞ�8[/�A��D�樉�$l�̐ۈ�m���r�~�����������6�nd�/u�z��߫Ȍ��6?�
A�['4��D'���e\�l�:`��܂�����Dl����|~p������D��[�l퀻rff]�ן
l-���s�`*�����uM���2��I'��$R	C`��d������֣7�_*`@�6GQ�e�!i4'_6��(d�֓96��;H���S��N.] $�	2'�@��4�18O�W�n��T�	0}XNB0_��@��]0�Id�n�`-�o0�`Q���+��J��U<<<��)H�Ŕ�uY[��fw�}��������R�Ep�D��).��}���,+)=D ��v>�b
m,�p�'kp&h�-�4�0G����S�hmW����>��]U�wb�eb�����K�Vפ���{��Z��ͼC^�H��"i�}�$�;t[Zc�u���<˨���ͣ�Tkzkw���'�{!D�-�ďS�ꪂ9��D{t����o�9�̊IΤ���[Xj��Nv�d����x�۷�]�ɷ�	L��K��GX߶�¢��r�M
��[@tM�,"�-��a۵?�!�R��Hd�yو�:WO��8[��0�/S���ъ�,�dE��T�*���YBrYllB�h�./o���Kt���ۣ�-���T9x���'~��i��:e�K,� `�0��0�tȞ7=��m�vo~����O��,쁙QUkc&�S��E��������=YHR�
���g�n�lgoP�w�[�@�ɲ�B�������Ê�%�(��6��=�k��jg�V�l��K����JY�H�{�pp���C���2�"m��a�?w>i�xq��D� �u�'UB���ձ�L)�|�W�Qgs+��+Ԛ�L7M�ə�yD��,��/-�fy��O�|��d5#[3h�D:��U������	��+m�@,(�ѫ�?q�O��y���E�30/ �������BWS�Kq�#�07fhfUQ[Aǟ빧��7Z=��Y~U����IԷgaA�x��w�9=���-��w���FD ·2��4��so����)B5�R����	�'�cӉk����3�<p-��|k�=_x#�Վ��7��Tٳ����j����o�ShT���@_$B���|�06&����Y���#���>	�t���0���n��>���O�6�Wa�0�-T<
�(��}gg�ӵ�C������H�%|��j�ɿW�P{���N��o�ה�<�;��u�}_�j�]]���{�:��l��ν���F�׮�ec>���mӢ�O"gy5K>�}�`�|L��	��0�s^q����^^K��LY����Zyj�]|�O�^�w��v1q��'k���y�Qo�v�s�n+K��МI� �DQugd�F�����"��oBh�9�M���UR;�j2.kԷ8E�;p#ր]�.T�j0��E ���}Y��'[�Q��P���A?�G%P���c!�{`�nwP��1�&���{t׈����)��E�/O^֏`�?&�>7M�ea�y���J?6\��[�e�2�,�H ��5�;]�����/_6�,��ڮ)J}���*'6��س���N>�����0%Lz4ʙW�O�ȵ�>��v��d�@?B"����4�|�uӏk���6�b�hw�$[@�y�}�g7M}v�,V�����tQNd��?�!�ct5�w'��ZX4�4On�45��ka���@�Z�#γü�á�~���Ey4҅a,Zn�xQ�6.WA��?��L�
�d�A$Ғhv�� �uO�3y��9���L����_��Ĳ��F����=��ҧg&-�03����K�ӎ��| +Jq)ۨ��
X�u����Ϟu�hV]���ă������1\�Wl��@�!v�)m���B�J) "vMu#Xq?����l�fFZT�;����)B�"�����)}$i!�!Ao �����7�l�R;�k6[ݠy�Y�8��VEV^z��i�����7�U�@L�ټ�� W��.p�:���p���J��K����]|�P
~��N;(x `�1�ۊ������6b�;;��S�Mr���N�p}b�%N	�M��	��	�&��b���78��n0��=�;i��"u.�����e� '�[lR�D�R�a�F�zr��9p�����ד��U?K����>��v�:,���B���{b@��m��,�?Z�\Sߑ52C���� �ʼAc�8�F8i{|�X�$�U��d�*Rx�\�cY�z˅�ADozcǼ~;{"j��Ʌ\�8s�����7�K_3�m�q�b ��syXOl��
��!t����`�����#ܚ�/:�~s�^�����6�������wM}�W���+�L�_ฟ�DK��I�ڝ�2�ǃ�nb�2��P�����嘆'�_8�~���*�G͆�FYȸr��Z���p׳ċ����٭��C�8�?�2D>ڷ��]i��V7�������U`*�Ɖ�b=�->X<c�ւ�ر����p%���ʷ�kPW��\���1v$)���wj���G�����yu��ـ\BЕS�(UM����b�Xzz�7Ooiؽ��!$_�n��@.�"�X�\x8|P�:^$H�Z�����w��� �;���
���\���R%CZ�`X��-�~��{eu1�F}�H/1��z&%G���uh�����b,ZF%�`�Ob<E�/�e=�J�����������Nͫ�;߂��ƞ��+�߃sUԽ��K��1e�v�����"A��D��L	���(�j*P�T���m��d��P�}r�YFY�#D��~\��)I�tFU��slF#�`��m�h�Hx�^�(ke_�"��g��o�WVĽ^.��0�"9��7� �-�H�Y���$�*â���{.(�M6��gv��2t_�3?'����DG@��ڸ�j���Ȕ�m���S�y�Y�O�շ1�D�ٸ�A\m�>�K=�� �/s�r�����/��j$ow��:���0��-
�,6�&I�+ �-ߦ��уԮ�? m
~�F'��� ��i�Di���Ĭk~�{�7��O��/� _��-��;��z)�fu�	����H;�9,��	�{����Y��.�����! +&�f#ؕ�����9�Z~�����2Hfd��_��L瞂�
k߀��(-�5��B����]ٗ^������$��n.���W����H�<�������?3/k?`	h�L�����Pey]�UN���N� ��vGO�c�p{��@^\gȻ���&�oU9ʮH>NIj���`"����j��΄��	kňj��ͲǼ�S��$� ��q���*T��oŶ�ZT�@e����S�蔄�cPh����vnET���J����9���VX�M��[�J/:�ՠ�J�w���!=���#*Z����ץ�.];Olf�7�!�l-�pC� Ġ\��C$���m��g�c���c�7K'ֺ��R=F)�PN����:}���O�,a�TvW�UN~�%�F�����{�p��:�My$�FI)f��p��w�-$!����ɧ}��̊�à���(���E�AF���N�ICc�3|��"-;4fC�G�a���s$�㺳�s3�|ͯxݶ�u[�A��܏���sւ��z�'��c�Ľ�]�d"�m�.�IRS��]����C���������^�.Wն�2)7�yp�L_c��A��_��ԇ���G��PB�?��پ�#��s�9�^���[͇U�6~�m�R'B	hJ|~0I��
{� 5�k�h���"��C�#拧'
>i~L�
��z�>ilM�?��+���I���h?�!���7S����R�6�'nK>4�IF/I�gݹfl%`:�f�T<�W��.�q�::r��"ϛ����PU~���P�W����9��3Ő���f7\U}��h&�x�S����N����v
�y��;�g^۠�,yl��`���ʸv�dK�s;�h���������K�Z�#_�=���I��|Ƅ�N�1�|uC�L�5��ҀH�@5"F�H��DZ�{���9��h��,V,�}]E�y:E��������7�y�'�WB������OZ2���˲3R��B�/o��W��|jǝ6�1��<Y5��.����m���P5Xt�����p/�{�d��TWs~[c3�I�"�lUM�����Y�B�99� �'�[������V:�q�`�\���08�A��Lr1 ���R��{���ueTٮd��a��w�Q�{�<�a�0�zq6�R���ն�=��֊��PM+,��&QE)A��L���][l7g^�4�O�qC�ダ���*�ߥ�������n�V��A���Ő��ެ/�5D|a�_����L��8�m��$�x�d;�yh�]W�t��r�<A;��ߺ�ʧ"M����p��&W�݊����_
 ���G����a2�f(��-�2�z��t�f�.�_���r�4p��u4�/$Fo`z�S�U@��B���U�&ig�y4 P�n�_�u�Qc�W=n/9�h;�6��Ah��X1Ga��M��]�����^�)��kWH�Rl23YI�]��_�)�q�A�-�3��n4W�	O����z'}ї���FV@�]�F��1�Ms+ �<�����y���E.�&s�{�b4���p����x�����n��ǰ��A���5��oY�@�O�/-[vP�tҧZEt~�-F�3�Yz���@����_݊֩���Nt8rK���s-92)j��.�������%���<4����j)7B�k�\w�o�y)EQ�S��o/b�4����fYT��k��E:�IY58\�����|Jn����`M�G�������2�(Mb�ț�G|���F0�ϳX)u��_���
��;�;:�oN��|N�R�6K����w�ܤ���=V ��s"#S���hm?�~�B�c���s-�M
�0X�A	Y�F�#�6�I�T^s~��N���$�}� ��e�Q�%
�߈���}
���0&]l��_��o�ѯ��1�* �1b�X��u%ō���90���?Rwf#)��S%ʔFbڡ'�Fm~�==fb�0��PMᯡ�'㷹��H��F�IE�탓|�fw�[�>X�[ۼK&��`�
Y������۵y���
SMq��v��eo]��=qPw�{��Ğ<>.��/
Rf�v��vms�����*�%ƥF|el0\_�X+��-��Z����:꥝�˸�E���f˾@�7�%ˬ������h
F�U�D��\��^����l�`Q�l���%u���lAۦ��F����}�>��~�;KL8������ oto�*}��-���@��A�vm��m���}玏���w���n�K��)	x/Pëg�u�q������hB�����b��w��*y�\�ٟ��)(3!չfSƄ�u:�j"�� h�?��W(x�|uz���w����C'�)B�``oݺWc��X���߳��<���������P�
���=��/_~���F�]�[�CiV[j/��u\�{��3X�bd��.cP�R3bM��V��K�6�l&�>W.�a���wj�1�ֲ�����LP���f�vt��{(���aHr(_��Z,�9'E؝j̀��і~k��t�+�89��*Z֙~� ��͌@��Xo0��E��X_�������D'ڼ9��c�
C���ˮ��M�ޫr� �C'y�M�1����i������f�	�����7&0��{p3�L�)5a�wu�g����3H	�!��?gҘ(�q`�R�ɇ�5�27|���)Z��P�bp�&4'�V����C�x�/�5��lX��gS�`W���Lz��
6��bQ �4�z�T�����@,��TLg����[�z�PD��%D�%f����ڵ瘀n0\+g��<c�l�������%�7�~N��A(351d���.���)Ӂl��DaA�/����Oy�2��1ƾ,i��2*�s�W.KW;%3x���0ơҽ���A�%�O���TdG6Xs��X�H�,,���ڂh���v+�!��l��e&�%X��~�_��� ������>�5���om����n�%4Ja�P���R##d�6�jG�"*�$��q��?�~F�a�=��wB��X����GK�(������j{��e+�:��xV$��i��R_���w�]2 ;�d����;d���\���[�]�u#.�m����>��ʇ�I�PQ���5{�[T���=i^�KٕP��W*@c�:���mU]6�}�ۮc�i!�W!��lB��C�3=������ǒ��O%�����m�vL�ؑlWG����7S��^����3����)|�Yh9�c��$���[�&P-�u;ݺ�7�R.��E9�@N�� ��L̃3ϧKU�:�����3���N�a5�'�"(�e����OL�����H:>Ó~��[[��f�Uٷ��7��H�Ѐ�G�<���▙�Q6u����p��2�'u8��1�;�����f��e;��p٧$7�hv(ӈ�X��^1��?��:-,��"*U���Y�u�ܐ���fm�Et���}@�T�U	��|*~Y�A$,s����lGf��t�j�u�~��\I���Kt��-En�:�'��\�����c����m��J��ã���wM�u>�]�2(J���䜷��4)�u?���EZW3�]���W������_t���eQT����������}���c��ټ�uؾ×w?��#��j��;<\��({����l|]�����/��a�*w�^�ႇW`�H{�1�4_��0 b	�?V���I��#O�u���}��F7��^ui�����
8�T������hIy��Ke�mQt�_/P1���Q�;���j���K����}�n��X cCㄮ;�(��)D��cSr���%r�)�	S��S*Q�mMd<�����׹q8���q�r�6xx�]��z�A�����7���8
Z�������[k(��_��W�k~b�f��+�,>�2�hWU��_h������E'u���Ht��u�2����7n����y�Hf����Hbݶ_#�F0�o~�}��i'���~`Ct@[�Y<R}���o��u�����2��	o��䩔���+�qjޮ���X��๶9CjLk�3v$��L�s���fWYy��<M�oT��n�I�6V���m�nş�	qMvS(��g{.P�/��Q���?��#�%zN�K�����!y=K��q>��1�<���}:}QR��X����ѷ�����I`b�_�"h�"MW�JX�8#fd&�o[�M'L�bR>��EQr��w�B�,��r3ʁ��ugv��^�)��:�b|ڗ�Z��'�@�1t#;aF���ê`^��P�D�����8�l�2�]HqWa�ňQ��h*�� Wzm<��<yd�
���S9XKɕ^P � ������C�Q�����`4[0 e�o�hj�n9R������v�Q�"���8��}�auT=;wd�_@GM~��W�3���^����<�}G�%�מ��YO;V)Nj� �����AqPڥ��^�%��9�3.)3`MH�������A�r_(Ťy��-c����������K��bN��� ��� �Ή�XG����g�垉��=IJ�:�D��r�� #���1����<<�������2 B��_D�9y��+x��CG�9���X���͝ɲ�<���_���ۻ�C>sb�P�9�bp��j�'f��Q����Ic^�z�����{0��Χ8�fU��҄7ߧُ^.�~p��\=�~�3�O)t|$��FMDfV�!yn�M_��P��C�'���w�x���u�k����(ll:�@^o�z���O��6Ul���)�g��W׺d��h@\�"�@��@d�{F�\�~�h�z�`��(8����@n�~�Q���M����G�q�\�JBr���C���~*�?+�� �uW��g~p�&�sh��_Z,�`������K�W�h��C�՜�|��;��ěg܁+��jQEU��r�Y������^j�<>�2���݈��~h
I�V&� "SRE�g�%��Gm���a���Q~�0���+�!�����K� y艡�$�YG3�P�{��>tdGSC�p�;)7�;iGE������5{50�@��7��hG�_����{���!������1W��w���>�|н�&RWJd	eJM���d�?��K T9'Ņ���-�O�*x� <�-ҽ�+"��s�A.q{��r�{M�-P�	�O�y0�I�u���i�=IL�}v򢎲���	���Ɨ/�P�!�@!�?[�M㹙l#}>�`U�~�$�Lqw�G�IS��] �Spg)���A�c۴��p�@$xB�����ht1U��:@�����#�*����g��y���k�DB�+�l�kx
C�T>cqܰ�Sd��:�eB�v�i���Ƙ���O�ȟM����3��ڷ�!���J�q-&[�[��Г9��TE���i��* ���D�{T���ն#�ҕ[�@<���n�*�8��s�m�����B�2�pD�S��C�lf��a9�,�P}���C�0(E��:��ˌ���C���5��Fe����&�_z�R�e#�%�I�ք*�v�+$�S�7e��ۘgs�[lvsD�i\��6���{OO���5�\!@�Q�T-��<�7-*��n�<<���Ud�g�����)̀�V�,�P��|{>�I�f)�(��ϟK;������B��<}�1<�9���D<|�0�ؔ�'�&�1��0^(��?��.Q3��˩ӂx��=zh�2���4?&��aL��P�?�PQ��o��`�l�L���D�A �[�=D ,K�,��Ds���>@�ޣ�`R�����8Ƚ���t�=;����\�R 	�"�F���EA����<�zLY��G!#a\��
O���j�=�Ӻ~���k��~�ШΘ[a���z�OU-�jY�;${y�ѥ��1--��'_��X2)>9),�k�%�f��毷����]X�𱤫\��y�x!z��l��
��b&�y�e���L8�l�Z4f���3�D�M� �E�҉��Y(�\"ͳOz��#��ۄxԻ�����Ӵ��C���,M���<UX5�%O�ڈ�lo��UU��%
T���7��������_�y�yPZ��$����o&�WvN�%�Q/�`��O
�����U����x�S}0�so�&8 n�R؛G��mz�oOSyND�7�|�a�4ko��`�����)R�ǰIˑH3=�p����R�����ת�xmm��� -Y����� P��>`�0q��0ڒ��xo;�V���զ;�i'Pg����ÈG���[1Fw��b������%���/��!O�q�*�o���u�
��+�$�F��tH�گ 1��X������?_T�'��`eR(�ebSq�g�Z�nF�y%邾�����C&x���kU�����ܣHM���9B���i��*.�*K��s�dЖ�\q�ڍL��W�����xa�w����L�����̯��R����N��������5��s�I�X!t��fU��2@�Cm��sN�џ��X��x�*KO�3� ��Vi9N��� X��BOa!>j|c"�}&��if����5b�C6��j�ɑ���=%q1#6�˲�Ȉ�S2M5��H��8���	��?�AD���u���'�,t�&��`Y����}�:���R �W������q�<�eeG���R3�����l:���$��$ٟJ0`'�����	&�0=�ⳋ4{�@�d����&�u���.�-�/Gz��K#.�rh��",��'��Roa��?�0`+x�@�w��&��r����;D�h7�Ę�����{�I�����k��Vb����%�ט[M��7$�k7\�����A�	h ��D��F��.b�#�gu@��Gx�<PC{>uxK\�-ፎ�*�k���;އ���]+0��^��8��,�`;X�qi\��/�Q�̶
aRa�X����㍆47�Ym*��H�KW,O�zY��4�˜�H��^g���A��<��)�����J*�Vs�}:t�т὘��e���L1I�D�1y>ܤGK�V���ϩ�2�OCP��2��y��h4�1��J	qīCf��D�Fv���`�a��	pX�} �U�q!�����LZB"�$�f��?��<�8k-9���S��9GҪ�Ԝ7̠��C��p��.���6Г������=�>�p��RQ��7�g�e�:?���|"w2��h&m<3`z�q���:�B��(��c|�w�Qu~R���F�7�L�[6�C�`���<~�0f�W�#h�iy��%<2�9��L-6�u��F�pa�h����M�] ֪������i��T� �z�� ���B�coV��Z���[U�k\ub��/�HrA�ӡ){QSt��ZfP<����T��1�{�����`�/5K�<�G��"�]����,��s�c8�'�\N�pRu-�x�6�����Cc�O(�e��/ŏ8��ZD��V_ߑUD�2��E���".���$N�A�t�j�)Y �_���՝/�&�+����S	٢����g�TE`Hv's�w�c��@���K.� �M�9�Z�T	�(��g�Re������!����6
�?+'g\�d�G�par�y��T�Uz���ɚ\�T��l�Hh�h�}0�쥝��ěol��+�v}�-��rz��6={顗ƈ�+���R���!����+��}u"+�Z4�<+SV���ό��7��eI��߮hg5{ϞJ���	ZҰ�跪Ȥ�� �ݡ7����;�-��?+jɌ;�������	'\8�Y�����5%��7o�.t�~2Mp�a��mB������nd
�F����c		\|]�y�jn��&}(�6�~���O�9�H ,����5V	b/q����$��9Č'���(9�E-�;3�+n¢J4��2�q[���&�#�YˌS�/_*��Y�aø�s�����i�[rF5�[[9L����@<�y��VZ6Z(P�M|)��L��*g7�2�2�WD��̐���8����Y���#����+��M.|��+�Ay���;����X�faE�o'^=�S��(�$�Z����B���>Ξ9��v����Ih����f�w�rS�3��[�2��` UUǢ>��GB\�m�zx����L�7l@f9��"M��_=�
hv�1Lr[��6  xt���7C��^݈�\b� E�Aj�4��ʨsy����.�S�z�8��oZ��Q����������#O����a}��~�o!����׺5$��Gb�K�����hk!���]�������� I���:��H�W�B��K^����>�eO����?�DKI��y�?I�m��x��� g�@'}I�	l����闁�H{�9�[^�<��V�5�c�C�T�����5/�Xi�3c�WU>�~��u�����[�����IE��I73��ZS�G�w/�+�i�y��u�p�"�E�N56�2��#�}�4 ��-�J��Ɵ~	{;��^>��X�?@��!_���|��@��B4�w�-�'�cm���B���+��HI��wD5:�.��
���7I�!Ϊ!N�Xԫ3�t��Xf�͖}�d��Xz��KHX��|Oˬ�� ��D	AHz������t?θ�ߣ�>h�\��A��<a'C(<A:ݏ����'	��	aj=���Q�N�~y�|`��'�-ޢ	��5�^���6�@���&U�ϕ]��JG�O<ѶwV��L�$8�����Q�ڂ������`g� '}	����̃krI}yH���i�Q�C�g\��27؏;ռ,�{oY �P/�������$���Q��1O�M*�*fi��7I_���Š�1(� g���-�!�;��ǻ7K���~��6�������|�c����m��B�� '
�~n��X��O����w��H��;�9 �'+�=>�y�+�'�d��0��`\�U�3���>v��#�õ�|��3f&��~��	�6��t����(����rT]Y����Q���O�ʁ1p�Z,�r8��t?ٸ��*A�D�G��/���S��!N��W��y����Z�����|̝���,i�x��W�a��h2��4=��߿?��ś���`0!����]�9;!�-���iC�J,M�MY�}����a�gk20C�������:���: �RvFH��:��eD�*�|��N�zV�dpP�I�,(�P�xKs�Sf%y�?I��-0=�"�!��4U�=u��w闥�ܣ��/���:;��	�Q�� ƫ!���U�V���e�Ɵ
��O󉦸��:��j�AS/(-���rJd�ui�c��>��Ԣ�IK�4;��	�;��j�zu�y���Nh���<�^��s�>] �������Yޞ6��V��D,{�$�"5
4@�~���p-�z(2�G�A�6�E^7re#
���)�ِ�6̹K1�O-�Hƫ94橇�����3{Z�@��޹@{⌵��]��.�2.��p>aҐ����aO��;��~�������̨6�~L��^2�*	�I��c DB#��Nb��^��(�j�\n�5Э�,�0n�S�qw����y5dǸ�/��GP'�W�&r��k��Լ�ϪE`/Aq�0 �_�'��c�Gu��:����'��%����r������8�u�br@���ׄ��@|/k��ƗRs�����)�;N!ۃ�x<��Q/_[�7��FB�@`�!W4������Mdm�Z���5���į��Җ��7�7Y(�99�(�= ҇���)3}�����y�vˑ��:��mN�觎����QT4��N;0�p�K�e�8-�m�Wf$�"�
�Z�K]E��/)Q������鰢I�_������P�W6��*%G�����Z0�������C��~����I��X��x3��tC���^�QCN�Eu^�_q���6�{��U"�2mxW-��og��p��750������ux	����O������Lwqeh�	��NT(����|���Y%��!��1&Ǫ����rp�t��m�=��/:&�\QXvg�AC�/��;����|��':�4�#�IT�i�J���w�0���f�N2>_��h1v�]�J¶�n�9M���{+	�[�#I/��c��X��a�4��$���c� [-�N�*������)B�Vf��Wn��aAg����֩O5. Eq��J.5��O����,'8�f��A)'ZX��U�	��
uƁX�F}�>�]��R�s��2w�7`�5�������/��>�ͣm4G7N	��$��x����w�`�e-��ܮ��<V2>��8]���f�vx���p��x��'ֶ�x�Ś�8���Q�9��w���i`>��iqH�/.���p8[�jVE1"�L����.�
U�(�O�B��u�����8��=�2][gb�����Xژ!?W�^jv~̰�;v�ŏ^�z9�''��-�sb2�[�;�VT��C�Ҙ���Bƚ��yq�MXU�u�����|(���ok�������y}b�Uv�׋�r�%�v�(_��eη�4�Ӷ��C��^4𕓬7\�D���r<r�,�p��Y<&��A�VS��V���]ay��wV�k۠��SI�?�l��3��	�5^��Z"����U^%��k4�/���q����q �}a}���%�ւ�߇�E�����ռ��c��v�S�M��|ׯ���9�`z�$2ѱs��|JJ�@0���K�H8�����|��#����x�OGó߮�G���4I���{��K�gX�?��~�1�_NmA��2�d�����c<�,-�x�7Qŀh/�}����u�A�y���)�K(���U0�V�#g�۪�ͧ�"�4�Gٯ`�����T��$+;��Z`S�Pw���		ko����Ys�<L��%X��ڗ� ����H�8ןA�
�/-���6�����oD@n�������7d�Lْ�ZJ��g�8� 6o%��ퟫ��fDq@2�KD�u�Q�]!0Fqz��x�Y �͓��f��I<|lw������_=��r���d��X�%�ق�r�Y�T�"<!�2���4�Q���������5�6�?�$�z�Ď\�ٮ, ����=������ ��T��u���5Ӥ���8`�fz���|�n���������7뀦��T�Ƥ��.�
��xsi���e���XB,�{R�t��5�o[���t�%h������I�cf��Fw���J��۲1P)�>�Y�X���Y�+� �.��m8��.��k$ߵ�����}�L�)�\��}{�����Qs�����J�(���I��׼��-��Пv�Ҫ��vPP8��Bv�`�Q��j^�!9P>B�6h�B )���%6gI��Ff8n����	�Ň�rii�����s���C�}�{��m\���K��+m��.�SB��L�ڵ�[��D����n��X6l���9��nO'����J�q1��\��F��CIy|~����)���4f��*衂�[��2��r�~u�|������;�ujy����Ǵ읕���/XDD����;U�+��_��n$�S���vv���T�����X"�O��鈬o�74�E_�V3����x66D�`���N�*��e�J���+1³7�dFe�O�K���Z��H��/�Ff��6��"�
j��\�*�bI �l>���o&����w��L�b��6�z>9�����00�#^�Kdґ��n_�:�ec�����ʲ��!�T���w��Q���]R��b����e?;�m�I(�������H��)�ikU�\�<)����t6x��l^T����0�u� 2B�G�_\�u�w	E�v�FD&�"�
Ƚ�H�V~�:�h<|�7���Bg�}S�L%fe��ܤ�L�p�_:�=#��J�x�&����ZL�ߌ'���B����W� E� 3*�ﭥz�M֛XQq� D
�7�r��0E�q����UJ����Z��<;OG!F��cVY��B&��f�n,N�B�ϣ��׳.��;����澸�7Y��v;�������O
M�L�^��)[e��1$����1�ra�G�i��*�])��Ns�2���e9:���C\�����ԅ=�+G2"w9r��F yUQ����p������?8�O�Hi؞�z*�_�b��&7���R~4�9O
(�_�� �L�!�6*�h�����h�g����?�ڶ J]�f����g�LO��v��{Si��@��OU����60DI�~H��\���I�u��^c�.�XM�L�$�qm��5w|�[m�6ak׸�R�}1����_Q{��������͌��2[y��-��J���&��f%[��b�N��7��R�N&I�.xH.E5� �����~�E�c�"*�ϩ����udcB�%B�U���Z�?�Z��5�Tj��4Ns8퉹��U�m(Qy�5,:��]��\lp���p�,gC0�amo�y��[ϰq�p��
/)g+􇙔��"�J֪%�gs�K��fKU�"���K�}�#�I������u�D]J��V�e���?�D�(�W9M�Q���Jq݄��vי	������\;��3>�Ə�
�w���U�G(��u���C����ׇ�V�r��(�e������0�3�B��AeU�|�g
E'��OL��_��F���=i\�ĝ$�[�hC�u�hM��KY�ڕui����J�Tie���V{�
�u)Bu%B�"�6~�U�:��r�|���}f��y�����m��Kk
�գ��B�~۾Գ!�fdk��4=��v"����9{�+��by�F}�l��x���C��.(��ܸ�
O�1ݚ������w�g�`�?+��Ƅ�����>�����bUb��!� ���QJ���[�q�Kb��[u��Vp#c�;z������+���W�����ͬ�S��_�±�"M�C��o������*0�sw� ���j�v�-����>yMg�n$��|⃸ti��S*i\��/���`��ڵ�=�����g�d1��]�˝��xU��&�MG��|�d�>�+}�ǃ���b�ya��̴5��%�˟�FR�n;E�#�v�3}��ݚJ��Lc5?��V�@�xP`����-<� �`WQ�x�S��xw�M��sA�FV��&�x;C �*�*�V׳9���p/\)��ƨ�)��#;���q�x��v��z�K�u�8�����I�u�׌����d$����z}�i��+{�ǁ��R{E~�F�5�@,�N4��i_�ǫ�о"�u|WR�dM�`�I���`$)�B�Ճ��t�\�^p�3y"+H�9τ��4�n�E���C������Upm�ѠQ��U����ifru$-���f�Y9o�g�,OKa��`����-��L[i�c���B�=�a����3�{6� ��p����+�r??,��=wh�z�c���L�Gf+u������A����zKP�C���A��Q��!��x��f�qX�5K�<���/o�0���85#�ԝ� �����S۞����8ɚ��u�-q��1h1Y����+$�c���V����^�d�E��Ñ�.�PI�!q�gԥ^����'�V'���#m*��NWC^��[��!��#F̙�;�w�$��mf@>�����y(���H�Q�U��*���Y�*�YԮ'L�t_q�yЯ^�,�Ɖ(��/�F���P��Q��3�m�䮹�o�}K

��*�uQ��2���+L��WN�A����0e���1�٬Z��"�cZ�n
J��g�R
�����F��B�����o�����\�XM��α�e�X;/��c��@���O8�ic��P���(�B��+;�ʗ�]7�T�u@*"oG��������s�\R^���̲-�8.��-L�GeT���R
�ˋ9Vs������Ŀ���:�d!�kJ�u��q�E0���.[�Y/��^/}��󮘾�R�ܓ��P�V�~u�?ö4��5A*���Ɍ�����<��Uhj�Y�;���*���)�c�X��1�U�����Z1g7�p��#�1��U:�C%�N��5�(�cȵ��񦰈?�ӭ�w�����������䵔.��p�h<��"(/u�(}��
G�g��T�[�I��H_��7�A��WlK���O��,*Vh_�Pih3}�7_�LM�t�hZĽo��)�-gI`��?O��W�Xf������^V���B����S��j�y,<5}�W ����'�Z��+�ψ@]KK��Ci�ۑZњM��/��*L�r�>���M S3�G����	����`d
��P�O�$��L� ���4�Ó�3�I@�.Α-S�2���i艶ͥ���F�T^Y�MtOL�+T#~�	�W�����!�P�;_�7��~���]��X���5p�"�>"��<�+����i �L_ظ�Bݬ2�v��ٳ�[�ޅ$�-��̬7���5X�~$�s�ʓ�C�����y���A�Fn�e��2����,JI6���.�
�t�Ø_�����0�5Zd��θ�����`����<�X�<�
PN�i�p_?�WK��~x��?�qO��7�P� �������oV��'��=�Ӯ��_����gDY��%�|��#��c� :sv�5���0�e7��F�%�|��kZ�)ʘ\�j}I;z��RvM� �eQi9�==�Ǌ�Zym�ˊ��g1gq�y@�3��c��t#�Ky� ��oٗ=0Mq�w�MY���ݩ��L9�"D�m�>3����[�~�8�,�M���^��Be=�	��'�~�8��F�D����}U��G�_�0>�(CJ�j�{�Ǯ��$��H�_)�V|����yo�,���ԩ�0fT��`J��w�	w�¹��u� ]:Q�뙏�ޛ�0�w��X�����|��k��	��%m�@��)�W��rnU�ӷ��¸��m��]���ev�8/��2��«ǰ����S�pK�
�q����f��>����%H!-G!�����/>��ok�M�xt�՝_�~K$j=(�PK   �n'Y�?HU!  B#  /   images/585092fd-6de4-462f-8499-92296fb2c536.png�U�S��]:��n���	i�F�;�F:�����n���n�x����	�;s�ܹ����=s�<��@lJl   TT���� $lL��m�����EA� ���o#��hB�]R���u�~�t�0q� xxx��8ڹ��|����l�y*A	 0�+ʂ5=�N�<5g��=k�K��"3c�����s�zhj>����v8�*����U�]635����D2a���Dc������M�P~��"z3����l�Μ�ws�+<����1v��2nh���0�*�� �dz�̗.�`;7)�G�fK{�"j�R��6G��e��o���<��Z��o5І�h��+u�8oi~�'�f;- C9p�]t���F�,��0^M1��D�K��7T��*��F&���Jb��{.����a���"�P�R�9)��H��G��3qx�N��
����=��Sp�IP���=YQ#��Q-��\F�A� /R}cЩs�@} 1���H%��4�k��(6K
w�Uxt��c��[?2
��Gh 6P_�-���(�QXA1��+6o����ws��p�&E�{�Y�X��"�UPӊr�K��=1��8��K�K o��H�hV����[9�p~S��}wuZC�p=3��GPZ�d��-��jn7��~�ʸ���O�֜�����3iZ]2nT�p�'/��g�}�iU*�k�u��V��gOaG���:p�r�N�@��^\��	^������N��ś���4��Q���S��g�S4O_��&�\k����ീ�A촱4��N��u3k&lE�&K��q!� C؁HsCY��ۆ�@�[<�I����|�h5�@w��6�:<��#�w�\�ն�iI�m��G������,�}�f�ԁq�cc}�zu���'�4�6@[�KW���<��T����4.IōˍY�*��1�ف�+���R	^��>�]Ư�;W��d���tV5��C�xłyx�^hE�윽���d���7��7�S�+tP2�]��1��E�9��j����60��Aʗ}�e��3�vi#�k�cNv���� M�U����D�@E���y�̴o�U�;�]�t��n(-�"�B�}�2v?e���}�;�{��'��{�A�/7J�3�f�#��{2���t7�0����-��'@~z������
 K[���ϗYSIܯ�K�>���@ �p�^��z�k�w}�}���f�,��sT�yzU͑6�3s�7G@k��1u���ˀ�k7��q�������������>տ^���� ݔƥC��,U:V��3]�u�������&C��j!���W�>ȹ���/be\~Ii
�l+�����`$E����Χ�"����O*������|䢤W����'mo����
��glFE��_$�)�xK�EC�~H"/לiVcƁ.��4��tFNX�/��Z�3���Tlڶ��đ�Q�"F�VV��ե<_Z��������X�>��ADr�_��-��2�M��[���Y�£����R�"����R����}�$�b�E��x�@#���H>g� B�ӆ�z��F�\��@tR�>��d���9�����8������N�1~��Յ�ly�H*�n(�d5��cؑLG�s3����j=m��� 0��R�ˋT�eM�-֨�B.u&o]��?,��aGYA��i�L�s�x!�5�7�������hpy*-�l�_�FӹaQB��s��c��ٍ��4?��\�uO��`�j�!�����|*����P�嵙�1�@m�º�t�:���g(�<g�3�=��u&?�[GG �ڗ���#�ڐ4�Я)ٯ.���wޅ����0����(-�A����yC�>[}5||���[�
}	~�6T�J���9��x�x�4DE�|��_.�1�.��l�6�Gtj��;o}B��@�����̛��/R��J�q
!3�j0���[@2���}8Cv��\�MV�iM�(�L���� �G/�~S�߳����������~"���
������ߋ5�yW�O�c�2|*��[���3j.-��ބ�"���rmʅ��m����߈dd��$NQP���f�546	{���|wRZ�I)/��Pάk$�3�6����~�RfU������u�ס��R��tT�6�u��S#����zd��y�w^�Y��E�'�����H`��i�1�"+�ˍW����	��W��0r䳒s~�tC��5�n�kZ:f-��j�7��g�q����7��#M|�<����
�梕ѭ����+�E}#
�̸sૃQ�z�� Q[o�伿��:!�ޗ�qꏳL���XY��p;~��~���ΩEMBD�sw�M�!-�j8�Y��dT��k���4	����c�*[��P�4�4�.����
�o���� ����x��t��������ye�o+w��T�g��}c�;�#<�H�<geζ�����_S��R��5pVSP��{���p��7�n��P��<)�ͷH:��uj�RAҦ�(�����ݳ��/eB=�g=v�	�U���62#]75Gd��nt|l��s+��hfn�ɥ�M�N�Om�"�aTF�'?֖旱.��|H"�ǚ����ϛ�>lس�r��L���޷7	!�`US=�>4�煖W�FNú��(q�asǟ�Tc��6P����Ie���1�S"��T.���n7u!�f4����os{kW����/w*�����.��%&�b>�p%�ݾ�%ߌ���W�'����q���O�Qf�B��!n8�sn
�~j~���|7�VU�Wj;CH��99��v��\QA���o�;�S�lj�٪V��Wf4��H2�8��د38�T����ėh#�f[����M@�E�'4�Yu޹�������e��7�e�ٞ�2v�+���?=��9)��Q�#�S=Bxo�k�0֔��2��l�M'}��B�r_�f��{�7~�W����<|KD��-C�4��Uʼ�jHa�
m����ث8��N\����ZS���Vڋ��G���瞾��l��zn����'��l;�W�m�K8G	���[��?�c>H���J0�c�����;�?��w�6g��2��(�1AQ���M�y���[�d��T@�i�-����X[X�B���f�0G�k�d�_��7w���1F<�l]�>�^��M�	��q����H�KzmY�82�#�s廛��E>.&�۳�ǥ�g0c&,h���6u*����U!��2J�|^Q����9:gr�x����]-�*o�F�̱�`��E�@�Jho1N�2[�^S���Zf�:?�t���T�Řl!\X�����
�0hP�"�w{ɭ��RiDc ;a8Ir���f�[��}�o"P�'��OG&$~��4��|nj�2��oǺ��Ye��!�<?��KY�:5�+f
���ɡ�8��\����L�����/
G�C��Բ�9%vJ������X������E���7VR/A*��sBN`L�p9#�(�9���c�J 9�O����FOY��a��k�IƘ�����BpBSLI�*׷�G&��gL�a��J� .�rǥ�6�.v�_mO{拃��~_�,�a��y6��@��4m�\6���B_�	L�𣖏���g�֜疸�TüO}�>�㇁���������>��	o<ƍ�������>�x3���H��Z;�)x��t���v��h䏲�Ws��ѣM�JgBSW׻/{=�6Y�/}�G�a�|Tၸ[3��9ހD�)l��?M�7�\ա��6���]fq�;�|�0@	�/L�IZS^|�a%��Vz�����9i���G���﷞�;5o��.p����7�X`GD`t>�-�Y���0��o���h�p3��r��;z�q�����B���^�����`�vH�%�%ͭv(x��X}�c;����}`����H��yL>0�`��m���[0g��W�� )Fr�Sf�$m[Kx��z�	�۫�G%�R�O��
J��+��F�]v4�9���;I����L���8��ҍ���wN)i1j���c�T&�M"l�"��L7�7���)=\� ����z�g�a��L*t�jB�g'�:2���������2Оt�raȧR��y����8��YP�Oh���a$6�!8n����,?��C'���.�M��#����nj� �~��K�nA�;�k�u�/@G�]S(�<k�lZ��Go��Ϊ��\c�e%�d��k�1i�"�5� ��=��t?���@��ƕ�8v���wE�Y������h*����r:Ɯ?�ms����l�Rx���~���o����~�F	�cں�?�Q�U
!t�����mEE�5qs��u���2�Y���-IJ���<��&�KC�B2���ʀ�]~*IQ�%.�Q>9w+3�@^�L]���`@X4���r�Æ{2�`)��<>nLʾ�Bk0<;���yK����ޘ�J5�A����n������HƗkh�K	�%,�û��Y�K�>�b����T�֓�P� � �ΨR�V���fM�{��;/q,T ���5m��'3��6s�׼o���a�֯b-x�#��}�q�Kv�7i�O��R?@Ӣp���/'e޺"�X��ɏ�����	-�*�p%����A���
�����?��nD��@�\�f�t���7n������XϘ��h_I�ˣ�1!^hf|�VS����.�'+�?߀>��^AP�fg��w��1!蘧qs�����xAp?�Ы�㽋��`z����6�'���f:�8��l@�
˺R��l�@<*���h7�Z���<Xy�{�#���L%�v'S~W��z��T9O���gc���k�U3�@�#���U�z����WAV����S��om�:Gx����U���xEf��b�J��:��,�D���������_��a��N�(����ο^^2l����j]�������#��Z,��^t�x��&x����%�A�9W�"�{~v}����t.�����H��$�h[o_#�fá�<�,��X?hr�x�IȮPJ�n�w�����d�&�(x��L�����K��^�BQ��lc-$����mog��v��>F���}�|�S}g(n�y,�\e��C}uv�i.u�����~Rm�*��MÀ[�9Va�/��T�ę�M��0�fz�ȁ�����E<��??��3�N�+fk%�5z
?�#f�(�*�����z��'�EH�
�:pơ���3tL-�?� ףg�Y	�h�wq3�wY��Ë�R\�d�{�����c{|���㄂<����/S��Y���f������,��C_�Y���Sm���ay��.cy`�n�͘����!Z*L݌����63�us3ˣ�c ��ݵ�h�~C%�A-�.�&��`Ƀi�U�H�*�~r,��i�'a����ӂ�����k,eFJ�`w�5o+���D|d�ɰ�KP��d�:M�`q��~���H�@K�y��@� �cidf�_�=c��`�b�yJ��-O�8k}��b}x@���Qr�bIi�\P3��,�a�!�_s�����K<����v�y;��j�WU�4 {��}N�b��&�$dL8�[c
������*�ܙ�8�B#F4�F$��*�~ᚾ>�IL��D\��7�6y�lHY�E��C)3%�᝶�nzl��ë&�G�$&Փ�B���'�`l *#��͙G��i�7dij�ߟ36�Fs��e
��xW�<Jj�i�y��꣰`\�H��b$����;�c�V��DRŷ	��\U��ͭ��y�آÚ,x�{��K��R?��E %�GU���:i�@Z�H�������٥�o�r������p��9m84!��9��q�P;���c������q�N���`�<�_m�_-�O�}�w\�N�Z6���ƾ�M��՞�������Dٙ�b/�BW�M�XT�8�y�����8CKі���8�h���T/\T
O�Z�V�L=��x���,��x�v����J%D�����i��[]^,��G�����>z�I1�E����'[�4kq����((fܒk�x�`�9�Ń�7⏑�Z/t1�$W���{�t��s���ܠ�UO�s"i���'�X3���>2�������O��j�#�]!���IhJ�D<]���������I�81��2��6�|q�iǂ<���Nr��;9w�=������8,�X�&p`	��9w\
VG.�8.q�EM�iY���@��q�1m�j߅6�}�	��Q��su��`�w�Q�i�[�l�!fg�>��m���wM$D^��+|>:��˖ޫ��Yߝ.6K�=0č�ө��e���h�s�{���x\��Y���*�f����\r.�
DQy:���[t(5�jM���d$���K� l#5�wǐ!��ɿ��Y��D*��;!��!9�wŲ)��
]�Q	�ֿ�/��q���������!H6���U�o>1��A*CP|�g����)v�J�������~A.-�rE�6.�(����$.���H�)�#t�U��+� �G����_��?���/�~��fO��)|rn~���S�Fo�7���R5��|���:�?N�d��b���g*-J�[�'ʺΝ�V���0��KӠ��K&H�'�������V����!��rC����ڳ˸��|5i�r$KȳA$��r�h�P�-T�'z�g��@�H`�;�<)�E�>��%^�H�6����n�����M���r�\�h}�*��V�4��Q�	����G������AR�M��G!N����v/0�����zy�����Q�!�WNqY
��o�04m�[�9�qQp��o�W�fSB(Ku��#�<'��'ϭ��gB�_0pA�bٝݪW�FX�l��I��N���2�&�?�����0(�P����=]D[�>302lv��̫��<⍌�^¤��q�Z�О���Jі�H�⿷~��[>�U�R lļ�R$y��!*�(ǻa@}Ne��`&<�!�I�ʐ���ć��m����+�&@�E'Hz9b�o&�R���&-�v�hyA��<�}B���Ҥg�(�!�%�jCP!G�jNnnD���ژd���.Π�i�U7L����\[���	.����!�A�{ Q�Y��?m��ak��f�1.00�S��!�sSA��f�%�Np��(�����-<��t�d ��0���	j�$L;j��
�\�p���ڱ�������{#8�x�ˌjN�TnU��f4��u�o�9�uD����F<R��e~�>�Kb���$3���D��x�漹��h��x4��a@������_Fc-�(��7���O h?��~I+6�~��/���h�Y�i��_�A	�������eT�$Ўl�U�3:
U:�P��W�6=��8K�V��7yѰ�*��$C�O�d�J�D-��M�S>EKN�*%Y9*�B絥���*7'n�JI`�CFʄ�w�����	C�:�.WP��1%�3	�[�lC�V��G�;�h�Pd��]4G���P��l4�=@��2����?�#N��µ��F��!_�Sm�4����dY���+w��V�r;�Ovd=X�~ɠd�3(,�WtL�jG|��/�B>�Gi}%聖3�1�T`~�#$���I��a��AN�'���,|bHM�3�-�"_�_4��1|���P��8E����,�@J��X*[)<߁�2���r��B�¼#�a�=�%ە��A�Wߝݷ8�^F7�fz��R�b�M�n-�k�A��\t��_P՜~f�MG'�sg������Rn�7�Ѻ����"��6�5�;(���~A�nԹ�
���s��6ݑ�����Z&� ���c�I�y�?�l����ђA$�͟��9ȧ���f��cPUg��	(u�>#
㏾��	gA̡ɁX΄ZcX.砮���hT~Q�v�z#���ph��'7��Z��Y��Z"��Y���b��p��2�s����hS5/W���G�h
=�=ZY5'���4��3�����WY'�����,Cf����d�:���*���#�W%��W�x�s��_U�I�홗�����1\)�e�Er,s5�r��YH�H�q�1û��@2D�R6���
�6y`jWDA2+9���Kf�L��9l.LU��v.�@�����x����X��񪼗c��`2�(	�N/΁����΃B�,��F9S8m[����Jq[�07w,+��
zE>�M@}����V� K�ZspK�	�щ����M݈�D�-MiuQ�|g�9{ٝ��|�C�o�k�n��Xdy*@��*m�����R�g�1R-Ks���9�d��j=s1�m��x�sms�O�1��[��Te+!�A�PK   �n'Y=��� Ѿ /   images/732af9df-f9f3-48da-8e69-a852eebc5446.png켇;�m�?~�B����"��)$Yeg���޴��޳���{�y�6![F��|7����}�����8z:��}]�y��k���~��KP�P(B�{�(��r����������|�{��P(�O�_�/��J��K����J�F�NOlQNNNl�V�v�Ol٬m��W�(P��ci����	K�x�**�;��Na����3�u;b&%�s'��b�<���+,��Sr��������u`��:��ënl|���N�o^����'������>��c^c�m�7낶,3�G���jW��~���^��~(sy���� ���������>���}w�7C�i}{;*;��̈́���l��EFrS|~�﷥�D����|���]�#|�P��J���`���P����SR%f�Ts4H.^����o{���On'�2�m��=ٞudB���7'����꽱8�0|�?�o���F�%���Xa��P����=}_l�������=�aq�%�A��g6�I�n�ו<I�����lL�ǕM^$cQ�h	g�i
�N�z�n�hP�K;�sϴ����ZO��Z��W�yVe�W4�m?hպ?Bj|���7!��\������W孾49Nʇ�/�xl�%_[[��������	�ʖ��I:q�3�"7��W����O���:�����]�_6�a�	�J�}}�.�]�'�in�H��?Z�5񂄂�9�Q.,"��S�܋Vj�����/1X(Ԅ��H���Sl��W�����r6);H���h�}�gR�T�m���IX�s�8�iq��������h�^W͎��֭r�q�dQ�����?k':�&G�w{�G����\P.�U��f$�>ނ�C�
�:�˅ѣN�#<�2O���rf_��U�J8��Ktj�_�cG�Y��=H��uA�%%Kll,$N���{�Ҧ������O�Bd�<y�a��#�G�Hۣ�W_�!A����~}]W�t,���<���;��.:g���RH^V5wח�zR�+��{�jV�\��f���W2�ձQ�e�T��Ͳ�bӾ�A�e��e��ϯ����s���EyT��� h3�V�E\&�bI^G.J[���sfٱY6n���b'�2c����,�`᫷n��D=�{�G��������CF��y�����S�)#��,X��H�H`K/�r[�('�|�d��G�K�������"WyxT����V�3\��y�����ǖ��N<ϊ��{���)m oK	�#{�+Зr9Xo����=wr��w:=v��U��<|-���
����WRP	�vZ<�$9^΀����\�t	�.��L4��L&<�� ����AH0	�qWRdL�E,�0&�M�4��%�g��E���r׻�M��w��v���Pd�a�k��Cؽ���[�>���|f��dtN(A����٢.�p��ݻ��$VǄw�g�g�W!���&^�BQ�2b�r��:Mz��
�~HM!p�j���7d_����t��,�<96Bں���f+�;}�6�rҋ�2�`��]�j��L���r^�2�Y�����2kv���q���HT��V9E���^a9�Q:�#x�e����?�b��1��s������g��Ь,�趽Zd�E�QZ���ut",36̥��ې^3�I����>�h6mf�� �1��jg�������racdCP������͛���,3%?��⃚���+�CΪapg%##vv#ڑ�?0�<11�{��BCƙ��@]_�5CEF�p��x�9=&I�O
�� ��P>>�%�߫VkYlh_�$�=�e�.e�y:%�l�L
���+WN�˧�}�3#��E��ӧ9����prl����	�߰���n'�@F��Z�M|J��o�+σ̠Y�Xh�{�D��w���HLS�%��9��n)W�
a+�A��Q���}0�7$�dTT7���#�h��&F|����E�>Nt�6{�O5|7�]�M�Y��q�6��&C�t�6l����Iܽ�B'~��SiB�Xf���'U� �Ϋ�̯�b��Z��S��Z�][R[Y��0������n�ըA[k�%��9�E�l���!��*&�2��ds��[�I�����~����t���)��&���I��O&��u��2t~0h	��hc���ѿL��<bt�ɇ�o�|�Ө��c�*��	�SesrY�9H�L�j�v�b9�I��+��M�}|�܅���Tl��X�`RH:��ߕ,����G�z���IG2ZZ�/��N���,yZa����<�2d��)�
�m ,8��Y�f�\R�v�u\��P2��鐡P!�'����e?/���P#dH#��#pOH^^���D��s�WYXd&6�1�﬌S�<��Œ��p��xr�P��mvg�p:WC�hB��l|ߐ�!�����XEDD��>H�>�v.�uM���Tb,�8֦*�kC��ݻ>|�������G�M�=~ׅ�l+�SPO�#΅����FJ�9qHB6�j�;+-5%f��R����}Nw$	k"���҂=�J�D}�J�Ƶ�ƣB��8�/;��5ɀia�C�H}��Rg����_��:tp�����kFo�JЩ�Yj]/#�9�?]A���A�u.2��|a���������ջ���7�<o��U�Hh���)�j��e�q8�F��W�SM���˟�+	���P��P���8$����nar���N�<ss2k{��QW��V/x�l���g���C��}^��#%^�����f�x�Ǿ��f�n�$1�J��'������V��k_8�n ��D��0��t8�T��ų��|�E>���u4���s�\��7��FJ̙�F��k/�SNnc����]K�?�����P�ז�A���c�`������'�n�44�\�i�m��쬭�A)0���oD�i��K�5'g_v�|��uN������U���8(�i�_�i�/N>"DT�XD�F����;�hf叏��O���WI�.��챿�0�KbU�ÒW}E�p3\h��ɠ:!%�UxB=a�~+�5ORLa��Һ�'Eʰ罤b��tU�d��xxm�od�Q�
�/�j��t+����:s�X�%����:)	���u�?�d"�U�(����U� Qv�}Y����+���\��y!y��-���*l&�����kW@��Ox���_�T��Arο��p�_``����=3��z.Ln��vY��,&Aσ�3\�.�P���[f~��b���	))(2'NDI�==��� !�+� {� F�Pp��������\�̝;�߮�`�ze�+@���`F?.J��W��o�,��̌�"��g&�ڼ�[k�R�ő4T�)�)+��Hph��1��$�>1���ǀ���W�N3)�<�"^�һɫ�6���CLW�J T�~�<a���v�4�/��Z�֊�`��G:���UM}!U���qW�I	��)[!!-ǥ!�q����k�:/1^ǇD�}���uV�އ�B��{�����b^����Sm4�����rު+�8OCr ��iEk}}�姺�Hd������B6�u&>�ܗ"E��
��!Y~X��Iܗ�A�a
a�٬�Z`i�2�{Kozz�TH���P�kB��dd�<���_�y{�F��g��#߾}+��0q�|U��J։�|�Ng���kv�����fPīQ��O���:��pT�s�G��7���>���y�>����&��^���S��D������\����1�F��o|[�NN�Wu]@o~�������{S�q]rX���~n��=Ʈױh8����«s4�oV@�"���p?>�pdp���}R�:��B ����`�������P9?@�p 9{T���w�f����D$�.j����>J�wY�,v%
�dS"�����N�>c��a�4��2޶r��C)�fr�*x":)�*��pnvsy)[KCc�z�qgNWL0]+�	����bb��*��8��������W�cL���d�*6-s���,M!��x�9�7�7���*d�r�ʳ�%9=���_r�Ϙ�T�
&�p���T�B�8
���A:���j4�d���������=�Ο|�t;�N����{�l���'<Ct���B	]��>���t�<7� 06Fq�m���s߹8�VW���_�N�2�a����'&��׈�9�W�Ow�W8�O!��OD���eN�ůZ�[	��<�b�*�%��=��,ڒ�IIHfzSe��v\d|
s��J����{��;�	�[��x��5Aq�4�p�(���Ra^��J����2.L��x>4��~])�9斾l��,��W���'�撽�P����4I��A�?�eL�aK��˸l6w&=��
���� &V'.������zVo���)k��v�NfF�'����>�>/��|�]�Y�Ca2��J�e�/�Ξ�{�Ţ�����-�?!,"2&;U� p��\���ca��.[�Ng"�6���ב��/-�u�o�Y=>��9"��M׍N���+i&UZ_l4�:|���0�ٶh^�.�!K��k�S���b��6t�I�TO4�*:�Ū��땶[�Ԯ�8��z��,p��1��:�Ji�y�I/^��6�}ڡ\�����L��e���q�{�m��.1�N�{zgB���x�ƪU~Sቃ�-pl��	:-�%���x���J@��{E�p���n*���	�6�ع�k��|0�?�{��}Y����lO��m�
�u��lV�9�\b���;11v�L֖Y��x��gr�r�aT���V��ק.���M^e*4�g��\Ql=.Rz�P% �ݖӖDmM��`N�l��wܝ�po��n���U�r�۰���Sj�@����é���|�$   �I�U���y����XM���6C]�\�s��P� �>�5��}P%�cC%����\��`������>�Ep�Y�|~߆tS��b��X'ƪ]z����XT���N�Vk�ʅ�7�1���;�m��wf�WM�(� ����h�KE��8��Q!�III��Z��}Zj 4�O-��W�w{�D�KEy9_�u�+},�	��7�>������w����]�����5{��i��q}�v��
(�k)R�<�ɻ;u�r�LMM9ܶ-�]7?Ҋ)�-a*��\\G�w*^g��x'�V��Y��޼:n��WL����5��8����Sa��a�����/��1�]]��㷱�[��+G}
�-~�L&,��!2�+�����Na��J�m�.ϭ�����:v�;�b�{�zbf���ˮ���:�u\�� /���@3K�!���^#44���Z�8"�����4D[pB9S�e��3��x��B�wE0��N�����aU��r��lR~[!���6K	�YY-eVU��po�b_~+l�UIx��_��>ҽ�����+v��fs��Hꩫ�W��
 /R%�H���MX7��m�-��D�<f���6+�x����=pX�e����Z$��C�m���\�F<i�V�"�X��&�}F�y�>�򛬿-/#x�|H������+D3�˖��3Z��.#�
(2�t��m�M���냜���~��:�ޗ���w@� �-����-�g3��hx�Zl������ƶ�i>W�S��r9��#��iT�����6ںmi�H��5�n�ieXb�����/^�� ܵ-?��4>��������Q�$!�!�WϽ3�1���
�6ֲ�fN�������K����2��7.5d�]*�j���OUEx���tS0y���m�CmȂ�7��<����a}8��w�4d�_�|ihkk�������CP�DU�в���,�<+[��#�᪎]DUL��q/]S�}��C,]"�o�/����g�����-��d֝(��Wd>�������q'U�fY�x��xm���@G��?��� t\R�e%�X;��N�j�����V9����?U�u�b��,�����L}FJ��w�\�̃vEF��HaD�zl��g���Fъ�xq���#��b6�V�B2���Jd[4����R|��AF��|퐱�AԂ�������0��@���D"�J/u���J
Hr�;88��-;P�ƾ7W��}`��TZ���k%҉<��"��f��TU���/e�y:��L�[��Ȩuok���ٕ�}+P؇3L��8s��w��9�+����98<���_&�}���p[�	���E�:"�E�Ĭ�,֑�Q��Qf������qB�Kbz���8K3���,�`�B�E��Z�*����]�t�j��E��~���w�3�ǿ|��p�}|p��`;�񅉼ysƪ�}�U������H1�s6xV�Z���34J���B�\/�a��·�l^����zeGd'Ԏ�Au,�q+��u��ߙd��dmO���쑢�=RGx1�wʗ��f�t����
!wu.���E[�ž�w�`��%�\�Y�}��T�'�R�Ћgg�WV���-"���kŦ]y�s��<�Bҍs���93B��9�.��Ta�6Q;���'={C�f	�a:O��<����Jj�Gu����@;�h0�_"�0Hj,[�^R

f��O���"�uǴ4�m�vH��
����t�ů\gu���k���m���i->A�[����6��Q&��]��c!���h�D\`e������pz��wy�%a�a�ؘ�F����&x�X\\�l�a{]0 �B�{��6��얃T�_]��<&���s�Ӳ�𤜗
����m��!_� ��}�*����!a�T��4%��|Pݝzj+���j�	�W����U���Ɲ1o�D����R��l����n,'py8#]��〦����h���c0�ŋ׊�:8�>#��Η%
������2ԫۺ�{�S|2揖���#�W'çB"��?�'��ʾ��:4�-C�q�sw���{�,b�u�:���ՒE<fwƣ�k��;	��$Q��QUMf ^��=�c;�^�������J��q<��(�L.#�ޏ)ɬZ�;1|�����XZ���B�`���e]|9��o
jAR�If�2�D��z�		��1%���������ϧٛ�M��8����Vu�������Ȓx"No2�ҢGEF$����m�)`_�T0�H�)e�ps尢��޺`�O)*�Q���� �ʲ?S4���ǟtȘ�CzR���K��d�`��\��F�ӧO?�� �? ��u��ڜ
��)~���h6m�r^���i�5��F0�B\U[����N$�B.��'���hF�JII����&ݗ��}-�K�����R
M����ܪWF��r4�52n���t^��%vg�V���ΨS�θ��v���"Ί�����	�l��W7V'۵k�	�Y:5�K�2X��|*wu����>g
 +K?P����E*��D��~�O���"�X�1���OƝؘ�k���;c?�eЃB!G�8!�����J$�ZT^��� ��G�a�@m��������r���d��d|B�H�����da�Ю�FU�7�������@��!T�^*r�u�(/$�,rz��p�~���!mc��ʕ$��2����l /˩�%}��F�����
Yj]	�}�� U`�ݽ��W�����}���KM-���N���Ld�K}�����?=���95)�eNv��C���$���ktNc.�3G�ѺHe�o���U������2�T@�׆&<W����]�}������*9	�q���j�ų��Y�K6008�����=v�o���z�7�8rr���4ҙbV;ƪQ���y�]�H+�c�БCC���A����~�(��~tt�]N��o>�}=�Y��tD9.r
ªS��tj߽{��h�t$������ &��g2ɩr17o#���K���iz�+��qO��?י8;��m�>�W�@������ɑp{E��V�q�ZS5'���F��pr8�f�Z{Se�9�@��C6��E	�E���¹st�9���� r_�ˬy%���\�Yfo��PF��b���̤�ԍ�G�z��R(�B�+~��bdؗߎy�[V�>_�iC�5��" �)�í�§�w#?�o�������<���dКZuu��pFeK<O�*�%@��C����/C��<��Ti;�L<��2g�����O�P_��DXr4J��-��SE�w�O���W�3�s����h�}ί��cn�Lށ_����}@��B$�b��%��˘
;�A�LQ�TT7�GJ�I��M��-�O��Ϯ]��6w�����ޕ�^3A��RԳ��פ���W��_a`h���Ub)�_H��Z���F˲Q#6���^�7o>�tXd�#��RSU�����74�s�䵲`.?��/|���pt�����P�u-G+U*�Vٜ0O}G�w���KH�<C+��}��n����Fn�n/����А\�t��9�6멬~4�L��<BMHä�I�V��i
�i..e���3�ٱߏZ����Q�3��t_�\����cp�4����0��������8/S%+�1�@
Њ۴��+g|��/t�YGK{����DP�����O"��|\�iU!	f�Դ-�<d���lZ!�N��A�C"�����_�KKKo|%Uh`��YG�Jg�9(��p�|�rW��cQkk��w/��m���w+�I7A$��_NU9����۷o�X��,�/��k��.��³A�Ӗ���(��1�U�7�u*yi 𐡈܇ٯ4�!G����<)$���kA.�LAH6��)d !pĎ�W9	�_�|�l������Ʉ��'���;����ZjV�%����E�'���ㅭ�X�Az� ��n�"F&��p\'���(V���Z���(���
Wb�$թ�n�5I&S�Q�f/D�����m�@���qgB(�GI�����&�hVٝ �$�����Ǝq~��sYF��Z ����H��8;��>�]]ef��r|��0_�!!�����;�+�,g�07���ݻ�*�H�*6t�O �9�>����{#@����̟��R6]�(6��N�?ޘ���U�LPR�;�Ⱦ0;K���pɤ����c�9�R�����r�G>5Q�KfN�P2�������7�4Y�zȹ��L��?B����_��(�P�v����?����=~�P(r5 ,���H�,U��@��𴨰�$�~G�:O�O��V����Uz�Ɏ����밤XI����K��\��_�@���.־]���֖U��3��WT��%3�r�4wd�ݓG�t�����j�*|+�h�t�n1��>�g�(��\�m~�N�[��r͢C+xJJJ�yS�����?�Z�1Z������4���7�o%rS����#��@�?�KB�KBOv�����<(G��_�T~�-C(|"��L�d�Q�*�W�H�.����O:�C� Zm�`�0�uuu�
R"ش5B��EpZ�����Y����B;�����w%%G�����:�����H3!����mN�u�f��ey�dӝ�����xXs�o��^�f�QP{�8>|�.�t&��:���R�];t�,�dir� �W=ˑ�*��ٽ7`��Ќ�+���qC�+?`�,*�D)�������=k��9a���O���?UDD�_t[����}:�؂����G
�p�l�|�ȗ*����"j��?KM!���Ĩ��'FF��@S�����D������4�/�/NO��tu�-g>v[��tc��5��I�u3�]*��V�
,֣�PPXXx��n2soi'##Í��T_�e6R�7[�b#sy��}0�$!ŷ����I����	~�Xo�4�F�����Pm��Bzr�+l_;"(��:ˬ�������S��K��UHG<o���Jr+�� <@�����6ip����	/E���� ��,5�23�d���he��V��rrt�n*VG2℧�'��}��DDl
�N��:��+�_�����[� \n쇶���͔�O��-���nɵ�h��Z�V�[����
�ڿ
�+�۷B���^���FӺ���{ѽy��װ�z��fs�=�n���������k�\��������D�A�����e�<Ӿ��*'��9�c@����(����r�ZQI�szz:X��u�]�d�?�n����.��->����֫������2�GG���B:�0��vLKxԍ_���ΚhF���%eo��t�ݘ���qw��կL�Y⾻�W�V��Ⱏ�(mq-_�vҽw�
�
&C��=r��e�E?br����p�v�e�ˬ��2VJ`�������yf�E��SȝN����t�_�B�b~~��ZX,&$�f�/<,l i-�8�`b�n^���,�:�]�E>*^[[�B&��0_ȠV�iA)�@�x��e�O`9���e���l3�G'$$xN~~�	qu�~�{������g�2�t��ϯ�����4$$�]�3�"�=��3�u��\���˔�Z5Ogt��bQ ���{	II�R=�z���z(��U�����փ��#'$/3�c���25-��6hn�iilZU���ϩ�e�)���)y��EGF�pĨd*g��=��|C�e�����Ϊ1�&4��ݶ���5$�D�6<c�l�	)�q��YY_���E���'��"�.��Z|���]�����%����8s�	�v�3�[
��b<w�d���Z�ץ�"c��J�,pmR�������Mh���9�0��L���u�V�n���a0�-9ec̿�(� ���@*���W��>y6
�1l���>q�Ly	�d0..�(9>*?9K�,T](%�
r�f^XSx�`��#F���UUK����'ì�[�>��r�_���6k����DԮ� (SZ�X5sLT�:j����W�V;�^��֠n�J&�%�J��G��hB�\����@��ϛ\�4
otCn������a����-��UQ8�]�ο0�`�x�j��P�L<!%���7�,BBաee;	��;�ޛ��vw�����q�۹#QO����+��w�xt|�v��{���=�_7� �s!yX�iڲ��#�K�3��(����XR���]$"�<��jk:�^}�lܳ
9VY)�#.nx�k}���럪e`�;(���M��r!�#�!Xh�5
��������ť
�9"]�@����7ϱɩ�S���i��'&&.�E��������Ua0$ɀ�G�a���	{��worQ����.Bၠ �p��qL��ܲ�^�Ӫ�㦐��������}<��=�tWʿ��t%��#>72,��Ç�Cǧ�Uu���G��m����2a=r�۞��kmʅ7��5K-�h���� ݦ�j�	elڕii�����zzzֱe^��?���(��,��۪		ٿvv_��E���靕W/p��2���������b#���ҲGټ��mV�\�9�C&$$�s���f��+�g�'�a��f�rf����.�c����}����C�Q4�o# �e���S�Og��=��Qm�ov�4j��505����{ll,���8�m��a���J��ާ��^Phc�sou\̲���������B�6ի'�8	+ I����)(����͉�I��X�*;�"""�&(���$�b����W��爣�[�ձgttt��لo�IaN6��%�Ղ�n��E���#�G9�P�#��������_���o�q�MSHf8(�u�f�F��C�U��{0��x@�;�'ܷ���@[�ЉWF�x��
ٖ����h⊹�S�e6y������D�ޑ|^M�:�N
���}��.6U
[���a���x�Bֻ�}!n��~\h=edW��%9OỬ7����f^�� ׬��=N�S�ُ�������=x�ҏ�����I���Ċ|�4�eos��t��U�|G��Ǹc���D��O��Z������r��yw[�{^#!����	��W>>�ѥ��"O��_E�]�:��g2@	�ţ��Z�[��9U.Ni1-"BMK+��R�WWkv�J^)��[s�\,���3�z�ڽ,�نI����F�k=�~7߮�)V���'���646zƄ��x�&H�e3�y\0:u?
�b�y|raa���ÎV��C�9���e�s6����W@���Q��Aghlh��+%�NR^��scrr2͘�a����tө�)���p�y�t����w������#{�fؿb@�+q�F:���\�9�����7�R1��� ����ZQ�w����(s�ώ�&�o�@�kj�5� L�<���e�E�������ȶ_�Mk�OOw�D@�~{i�9Z���]������w�!��ݻw�ϟ?w��1Q��3V���<��׻�!H3s���惹�������{ܶ�L��W�Xa#/h��r��B����#�11|60KQL+`|m���%�Oll�*7f�OЮ��ζ�� �F�+��wd�Xi<y�eyř <���B_:/���<MN+��@���s ����?vw�Y���. =�x�aq#kq�ow}��.���m��3���/󿳫����r[�h�����w��"��As�H�O�Tj�+Y���|�t����n���Q+J�{��<sK��*��%���.�!�!�/AY�0���;�)�t�1<xg�S�	�4z������ym�9�AƊꄔ������|��� �Ĭ�I( g����j����b�����X���� KApJL7G����v�\׭w�N���������s~��@�˸#��ٷ��[���.�Ͽ�s���<�NU��Y'5F�F1-?�vqƄ}�Lwd��1q��իW+!��pppb�	��B77�� DkhF�x�ܕtlv��Gnz�3����
xr�$��G��?o\�K�>>��h �E�l�R�(���GDD���刺�Z[Kt���e��L�o뗞>�*���2��I�����N<P���am��d�f�j_eb�u\"����\��/+�����C���LT��2��2����Lm�~�HSR�Ŕ�V�IJJ�L|z�����Ӭn�=<Z��I��ev����gA�F��,��5�#M���q�~����cW� �v�g���F���|�����WGFA�!��"��aq�vy����������|���}XЛ7��Tyd!���-·?���}/���Y������0M�q����~��?.m�m�[���O(2(�㷐��`V
�K��b��Q|vk��S�"?�Oe[[�=?R&#I))Q1�!A����������&.�ͩ)k%�-�PG����n>�?k#�e��^��]�	n ���2
@�]�GV����i1��dA�����3��)� �o�R��kcc+гAk�u�K֟_�#/���9���M�`��@�fg�����C,Z�C2�٥��t>E�coS��]g���p�{ȴ?S��t]��9B�(�����e����<�^�%u����A�$�${�^9�G���,��j����L$�V���ڎ~�%F��y?����F��j�N^���w�+W�������o=��{�x�ָ9��~���7 `0X,�B~rYY�p���ܓ,YYY~���|D�b�u��M�ࢻ�"o���y�$_�?s&\b"f@�`iJ& $��x��7��L;������T�`eqS���H5�^�Tq��������h<H���9�a�X�ijzZ�y��.�7 ��;���������3$�
!e��#�q�{0m��l��S��b G�G���n�ir�S�͈�f'�x��p�������y�@���h({ŗ�8�u��h�ûv[���`�zu�|$[�l����R ˹D�6(-����*Iƪ�-� �i��vv�@�5N�1�z1d�Ā��}mh��|ɐ��\��(���ubZ6Aǥp,���*�ɘ���7����Z�V�֪�P����Ň�T3��G��֫���фi�����Og���0'���'B��T#CCC@f�J�&�p-;kQ��K��,	b\�յ�{������"	t�	�*T`�PPr�l�L#C���-��F�����w\ ��o�-�xEo.*�|A^}�A���S��ɢ^t""�m�*YD�ԫ�j�z��j�UZĿ<IH�zy_��ꩍFn��|Ϳw]�2-D�r�@����`���j����MƬ<t����0��ȋ8o�E�v�t���k�C�H.���%��d�M!�afx��C��67�g���{}��ӯ[_��M�n��s�]l���ح�U������}W��k��6v����]����͑����t���ӧS�yN$��Ȱ=ڝC��?�aS�� H%'#s��5Z���l�bn�U �E	)�6i�ī����a.�n;+)�&��ׯ]��<��o4++KWA^�(18��ӿ�0�P��0���)�`oA�'ȩ8<���mk����ؙ���y_���Խ$�h�<44Կ���'nf�£�
�n��H���d���7�!�	�JH�i>���kll��̄��qgR���l�����B�'x�-P+VH��99��#>��Ȉ�L��܎�hN&٘�, ��o߾]*S�E�]�?�:S2�SD0�-�M���(�t�|:�TP��K�N�B�u,���𢶟aB���7����7�fdR���'�X�ߦr�����J�0.s������6���_�.2h�[�U��Op�.z�bfIYg��gY:��ѣG*������݁s@K�y���@2�~_�~mL�F����[�S��uw��ɞxM��dkk�od���=�V����7��<�!$"*�'N��t������
÷J:VV9�SK!]�)w�Ҝ����+	�f�?.���j"�Pn�D﵏���p[321P[���a�����p��o����e+�w�~kf��[��G����V��h���Q�$=�5󥏏���,�3����6�eo�¢"ZZ�&ii�U	I�W��HHH�˭����;J��*�<Y�|O
�?H�(��rk[�_��n�!�Dޡc�O����?�����,������������
@jvdw�άm���9�<�����AiZ>$(_FF%I����aU7 }�U�������8�f��d$�$(��_#�y�ӏ$��G�-$���o>�v?>܁Pv+"�_:p���U�=�Z.EϬT�^�3e1&�Mۙ{�y�Uy�ۛ ����t0Ve����g��S,_�`ie�h=R�0 rF���	R�2Mo(yE���!�-=��Mg��W��DS���� �_��b0��D��Ǘ]�	�Ȩ��j��t��֮��𨨨b��
�aaAg)/���/��hff���5�jkuV*�hUڛ�b�'����)��T�[���R�fg��l+ʅFk;�
���{�|%U� E]>2��4������746�Z�\����X���&?y��e���|J0�T�h���~[Fz�m�äm�A_�?�Qj&�����8!vq���Fr0�nڎ�+�n���O�a�⯀�3�j:�l��s�)0���������r���s�
�pH&� r\_h>�}���0ZU6$���c\+J�����Lt|��f��n?���Ǐ�so/���ֽ�<�5� �l��Myh��$�<�f��� !MB��ʢ�n��ҥ��=D^��A^����tL:�#���/��2�Z�oڿox�)�j����=X�e�;�����/6lA��Ce�v��� �g$  ��4jX�'����ϕ�^Ō�,���ׯK��;�`0Kc�O����dP��k��N7.ߓ��>{��eǛ�gͥ(,�!l��ރ�b����1;������Q���08:�-��Xx����?{�b���R,Ԛ������uu�ë�V�54����o��߸q�v�}@!E1BA�z' ��6��[���/P�x�5-�ob�1��WZ�<�x'�@g6�C N~��Ғoc0�n|\\esQ��qb6[����Ё�!��k���}�ρG�%�f�țc,�D.cl�Ǎ�ޮ��+�9�Q�h��IjMU�֣䷿�|]���C�]�������z���7/���	�8[H��A]/V�������lg?��9Ya�ק0��6`�B�hm%�~�����~J��>B���0��򴉚��gY�/׸+i`��P 9�����ɾƹs�~_d�\�>ON�$�s�\�P����h%u,?ţ�����_i7יGBBr�5�GB^����O������`�"l*����C�.??#��C�����I#v��;��Eoiݿ��R/�o"��1��ذ]���C�R��۝K���� ,��*��
Nr�,uE�9�C����N�1i��|*�D�x�7)�������R{�e�8������Gi:�9K�@�U��է.�0�jնw��"ͼ�C��3ϟ?��v~��ޮ�(c�t��#�ͳԣ��)�湀�]*"yY�-֔��������ڨJ���(F5�T.��&�UOP��RAm+�?U�e�%_��N����:^CC�*8E�(�k@���6�Ŧ}"
��B�g��O�E���˯��`j�כh)�W���:���R꜕o*w��_�j۫�u�n��gM������P���Sv�GN�<yz"Y�� �yc��[�t�_.l9��QW��>�mz�1&C��yg�������_&�ktQ�pڇ3Y 1>�����#���8w�ڻ�|���3�>��U�V��Ҟ�Gn�b���:借y���v'���*�i�ԗ9"\~�X�V�%B���S)R��W3ZV�mf��?�:�٪͞�~2��l��z��
FDMDDĶW�	yG=&f�N���͸ƛ�������GGG�y�x\�++���ٴ�>��*^+������8n�׬[ ��X��Ϝ<3�"�����zD(C����[	�öKM��[ '�ȫoh�? Iݰ��7��������	�q��u�._�t��~A1�ea
2�J/�L+1$���",\�d���ݝ���i���<2�[���(�����<u�4i�!F�MPp�k�4 ��U���ǣ�}Q��\%���~��"�ʨ�c��3III����*��ۥ%ض^G����E҆��.H�-��3-�-L��ب�L��N�c~��<�P����ҡ<A�O���^�4xt���Ul����w�n�Տ� "�cdqUy�0|��Gu��ˋ�g��:��$U�ɪYzOE%�S,��i���7%ˑb��\�BŒ�<ݺ�7&�sK�Vu\6{�Ǫ]�]���W�"������{$OL;�N�*��cOO?�	5������V��ꎿ��\ԏ���\t4Xw�py�ʍy"��!��ޡj�����e� v�1�k��A��3�^�����m�Q]-t��,��%��y��Ԗ�����~�W�����)�Y�W���KY^xKUO���� ���ү���j��陃�%7<<�J�(�Gw���O�F�E=�M0BJuJ͚�/?�؈��Y�F@IOO&C�n��J�v�����I�wB�˽�Yn�>�E�˾���b. O��7��;��
�?"�q�D�zԤ�a>�¹��ʡ��P&���yH��()*F���\&��:�k=z��_s	ˉR��Y��!"�b0W[S__ߋ	�a�D݄��g ({&�qq�-��Ѐ����QWgg�ƚZ���qںN���"��jx7����4/�������ݻ��yuG{�xg.�}l��'����҈�n������~Gr�c�H��.����k�+�����v	"" 9[z㤿�?�nr��I�յ2���W���o���!l��Ô@��������-�O�|U�ı��chdd�����bX��I�J�q��z�Q�&*�@��������S���R�K�*jjsC�v�ۢ��.�,�k����b�ҍ��g,r����>)()��q��H��EG3���yC�m�a��.���97ia'�:�θ<m�b�C�ϡ�Ò�D����!� THR��}��Lc��Ur�nKz?�	̚��>]���}�9�QHt�N�K|ҕ�\&�ؤN��U�i��d��(�T�<'�3��\�l
f�ֈ��(ﲀ?Ѽ��������Ut]�����"�!   �!���tH)Hw�
Ҡ�]��q(EZ	��!���H����</ܯ�����k���={�����ɯ�r�]\d{t�&_4���G`��z�w�p� �^�$4�T�求�Ӑ��I�r��Y���Tw(����<��������SR"��� ?�������SV�~�xq����?Ye9Z2���_=�t��y�_�qsK5p�p����:~㆛7	2������x$�����eў��S����j�fWW�ei�?�����>>>��W����ǁ��;5]ɫ��R>�t����%�H���a�d��J��|,'�@Tޑ/ ��<��Y�ى!h�z�u�x_�Ho�\�����,����G�@�w$$<v�8o�Q��'j��j�!�<�D���|5���W�����2ξ����a
���ؾN7j5�x� ��1�L�%͇+DI���o�r���U����b���0�����Q-W�:��E��M���
x�m��l��Uf��G��J�h�ݠ����l�$��x_YYݬRTU�X�z\�-���A��&?�SC�[��꨼�A*�^�?���ʑ���sѶ�Σ�<�tq�����6��n�g���p�d���|�˺|����,�y�;��v��Z�ƕp/���Q�'���Nv]7oތ��m �"i=Qub��[8�ov1Fv��w���E�8+�$q�C��\�\��ru���\�'�(�X��5�]�2)ĺ� �Zش���8C�G����II����o�����ȫ��V2$,,�I>V�­�;�;"�ң�����?y���͝f�����'�kS�ii��SyH���Ȗ� ���y 533'�Ofz��1��ܜ/(�B��&�x�b	rV�����@`�������f��B���p�4���W9�t+��VVT�;���Fm����k�,���$�ݢH])�}�S|k�[�r2���it� ��1C5�(�t�ɳ�/ۇ]'�넵���1�POuS��99�������k��/Դ��U~��6P�E2�����r�X$j���f��ٵ8~J�	E\�
�`mP%��E��|B��E;���[r/P�����V�SOoq��m�.��S�#Tt��e���w��IA��;�����g$��Q�C���),��ŞE��Č�16������A�=��I�_ ;�hh�;����s4j3+%w]n={�o	{���U{IABB�	�ȥ��鹡��~������<40�Bn�v*S���!��6�� �Ӿ?U�7��ļ�p�!� Bl���dPJA^^����X%(YI|����g�  ��O����aJ���r����%��^�G��ߴ�O���I��jYYY�yx!f8�����j�ϑJ��|	��>d Md�3�-�Ρl��M7Q������o�̒і��|�{���O�mZ��DE�P> M��CRf*�?a�| �s��1��=��`!�s=yt�;����w��g��j_�t�?
`#�NNN��Lr��ENٵ�~�����M�ؚr�Ň� ����3��ՖOt��s{Ӿ��y"�D�y����67�A1��ɯJ�}�p�����Q�s��j9)�b����gIs?��ګ��TH
� AX-#��(�6�QJP�AXI#� SR{�a>��7%�uc�)��$���]�uH?�����������B�mz�υ!�q�&��+���a�)��bV-�|r�QN�yYjФ�N���)*
F�{<K��h�̠OlK�3W>�+��j����G�J:���+0��[[���F$%&~}��s��(̮�*��u�*|��~�wh;N�+՗uh�˰�XN�^�h߷�ޭ�+�Rd��ݯ�E]�h�,��=�~M�u��k�r򋊬P��`���S����y&--�X<2&ww�
��#���-
���	ЏW۟�۹
P`��ذ��W_�t	`�Un�i@��TǄ4z�Vu��w�>��� ꡩŌ@�
���\G}Ƀ��u��Q4���f1��/�'j^���{�C�JJ}Ij9
�� ��s[YY��J�E�!~��E��#&+��v_�k�݀�m~V�d5�=i{{�A�Z���'/_��4����k���M�ư���w�l��e$X��C~~w�6���L���?���E�m�C��޳��`|u�a�D�E��%5�**��\�����F��_w�E���-,i(�)����҂�q; g�����4l?R/oﳧ`�����l�Uf�ᖢ.���v�J�@�Y0�Ł��>�Y� D��F�����0�K�d�&���r}�~e~[������͵'�Ty5�nt��

�|T�Xs����6����~�`1��qῑ�M3��������*��#���|#/�n��"\��DE'��|5惙�4�;3�@���7�=x࿾q@d'o���9� ���OEGǽP����J�o�D���jl���!L�J��q� 2��O��\`���;�������i�z������A?~Q�p��A��*�V�k��@_��[���*���?)��c�����uE�k&���G�z7�ߒ��T�c�u��{,�3���>eȜ	ݥ�g6:1��b��2����B��xT �)Gn�J����C�,�얓@��bWM���_HY� �g��%|�>���e.((���D���Ȳ����!���'פ���%}��Q
�5�}�T��&��(d�2-0s��WI�Kw\
����壀�nVkNëݘDh��\�(֯x��{o'hm�fi���GQRW�?��Y.���k鹽ĭvA�J����$��A�.w�zч�����B��{�@!�D��W�cl�4���������x��:�|8SW�/^�'��X��W�2�CI�[�2��iih8	ŷ����N3�,(X��>���P�:��"�I�L�Z3��% x��x�g��픘%��f"������W �.�νf�<��O23����$�ڲX�����sV��B����)l�`����R�i�!��̨�[�h�<��ls�#Z���`j�-Ծ��<%� �;���M�\+���5K��\
;j��d�u^�����,ߪ_L]�ju�=�W��jb��Sn8h��n�	�W�K�J��H�
�~N�$8�5�9�Bo2^�*Y*���w���;;i9}��/�?
#�PbP'L	�`Q=[�W�C!"t���6B��R*Iؑ���AA�E��N��'0�4���b����#�l��;%wµ�h������7�gU['���R٘YYY������й��vJ$׬?��N�������3�x��P�J��vF� <�{��h�=�F|���(���w���Ot����dǾ��rg�'�;�qqq�6�K[j:푀!��
�M�!�|ROB�����-,�l�K�:}��;��xO/#��Yر���۳2�Q���6f�,=#Lz
]�7S��������{o̚����(W�Sq��~��%�<�sy ���#��ȑ�z�B�1[�_�|,����S�ሆϟ�<��!h�F΅3]Jqk�s�;��2���Ov4&n?��Q¶T��KM�S ����A^�	ߵR]-Bdc���_c��*pcH��@�6'�5Rr��i��ӻ����?~�̩ ;�@O�.ؓ�E�a/���ю��tԼb0 ,�k�}�I�;旖�"�
�c7��4�|^�eXI#$�8[�Q��@pv2����������T
W�$r�l�̟�.8�-8`�߰�;Fو*��rJ�����{��p�������di]��_'�}�u��2ι�z8-��Jr2������.r�H"�gaY�&�'1:ک�\:Ƌ�.P�Zr���>ˏ[L��Ҷa9��h{�1�\:<�'�,`��}�SY� w£ɪ��DK�ݵ���x����
KkT1�H��XIn�nn��Y����>�ڱr��U	�0�`�|�Ɇn`��{W��F2�}�QeD�jE�ɐh���:���bCb�6UTȎ������� z�S澎��7��3fff~�	L�w ���BYk����uuu�gf�-P������f�D���8��N�/W��ܣ9�����_N(���ŭ�7�9����%���Ͽ:Z�7J�4�?�~��������#�3��{4�����~yy��i�Ǚ �4����o�����W<( 00�u��T�~�ښ�N�9L�vO����۹ �dv����T�w��:��'u���-�����l���6�9��l��5ȃ��H�l��S2J�� 4H���t�UQ��������Ytg�d�a��h�a���#e��'rrDjM{��Np��۬�rvK1��=E:�V�8 \��p�����ڟ3r��uJ�K�;C��`�_c�2�M� �[z�Rs$w [��H��ѧ���M~~~-���+!��L�ђj%�ZbL�e��.Q48 � O5 �^^������Ġ Ff�j�\�	�������i+��.$ٚ���h=a ��#,� � ��t�{x�&����>-Co&^�>���U�-�����B�*Fit1P�~%�J$��/�||U�er6��W Gt.]���SOf�'�a��b�����"��qP�^�~"�Z���`b^�� �/^����D����R�/aP����eu����@���j�e��d@��q�է����36΂4�O-��L||��(�Z�G�sd����!����1&�)�Y�L�<
$4��1_LML��]%�[w�V���dc�	
,����B:S����>�[��A����S�wv*��]#��W��_�K�c� d,֝'ᝁ�E����!�@�t^ib�e}��1�S�d`��E�<|�-U�����%X����v���1m����3��Nyx���Y�����<���,��$$@ ?54讽�CЫ#�=.%J�w�1�L`�q��?[|�X͂0<�� 3`-��Zh׭��Z�o/��Npg	=�M� ���p'2�����_��N=���<��|�n��u��=����3�m��-)i�A{	N���4'��EM�{�xW�	���#�}����(S�H1���R[@W#:6ݽ{��/T����ci�|�e��*|5b#[H�o��%�����.p�c����QΣ��RϚ
��kt_+�aw|^��-/W��%�mf����CBnT%�9>]/��������R���X�;#HD�#F����DRj���r��p��Q�Z�p�f�.k+_0�U��9*#��QN�f�!��ƃ�JB"_O���)*��˼҇��k���P�N�;|b�d��~��B 2�>�A�6�!�;f�}��qQ���(
�ݍ��f'm-�5>���Z���H��K��{y5b]����>��
��	�b���Dɾ��Ç���l7�����_\��:))syy��7!!!�kkk�X~�X������n�Д��>DG���&��3�*���k�'幔{��M`P���G�_hk=�8�����n�Qn9�Y��%�'�����3��:|�NSpE&�ax������(\0
Y`�o�k�z�Xۻ1�����GC0Թ�b�:Q���.���ղ*��|()�E2���_�~�/�*5�b��>�4�g0?7��6���=�s��hC����,��8`�2��ʎZ;�������)�3�IUJ2N�;�M�tPl&��kv����_��$��/m�����j��y�7fk,0����u"BB�G9����"��Qzi|\W��hF������EPPА�����J~�vW ��5��*h8�\D�x�{[L���,W1����<�F\~n�vP��(_2�`k��e,�Hu�6�7#}�E7�����^k�������F�[g��?��g:��L��9�gկY�܌�R�D���jo޼���z�u�l���ӧO�����
!!�P�2�8	�P�2N���Y�w,�(��^�x�����i�lAS���͕�}����_APY�޴�!��pn?;ހwX�jk�1O�[ Y��*fr��6n���_Jq.Hv�����"8��^)v���(X`c��bbb���.x'LX��ꛏ,S,�}OvF��{��_��[Yڰj8���6#�̀�
M���,�����߿	W5����N0��y+��y���X,�R԰��544���(ONv"�_hc�����fy�T�͕���2@V� �AT}2#��HHKKsV'Q��(���}�T��o���r`	��s���x���p���\��{px�Ɉ!\�𶩆|Vf�ೃ~ߞ�8~��Ơ������u�~1�ȯ��c�b�$��O�WW>�m:�)���=u;��"g�M�wn�,d�ۏ$�K�l��Q�눠�<q?C6(`��gV����� ſ�5�P(
d���`�Ȳ��>	�]�/~_Lƫ�==X�3�n7��*:�F<F���O���Z}�l$��CG�kL �\f��%=�,�}�Fl߯�t�@�cl�i�t�7�Q�Q}�1�<F�~��g����q�YFM��T�<|�a�!�N�Nju����§�����1�2�ޗ)o�Ј��t��~��j�>��{\��/)!J��������^��t�+�^E�U�rr�δ
֤B9��g�纑'��~
��H���Y�{��:�~���ǯŃJ����n�}c�)&��༚b�n���W=�����اA(�;���/��޿7Z_� �f�{z{��-Kc��;���j+�zKIAa���RV��'�;�w����"'�"��d�\.@�Y�rbb�)����o�tn��x�ܔ�*��"@�%� ��n�Ҧ�Dx��&8~����� �U��E�g\Zz��&4d���X�\��˪��P����.�lgd�5�u"���������A1&����mˤ��{�^�߀�ʕ�������!�b[saaa՘���B`��J������ì
X(��<����ȥ���".�w�~��m����E�w�,�#�����Г#���	>%4rpt,������̊��OG�)�5AN�U����>�\$Ί��N���$���fg;e��ꗀ���@���+�v�gP��$� n|o|�?ބ����D�և)�<kx��İk��#�>��;�3Q���Z��ϟ%���k����x���_C�@j���N	�����ʪP�N�~B�"G����R�/�:vv�����ި�(�e���w��s�����6}º�*�)�]e��pp�����<ū�#|�����,4 ��wrU�5����Q�	H�����ԑ���۴���>�C��"H-���h��4�3��So�����R�)&��7
˓��m:����F��+-u��+{l/�7�ou��2A�����hT�cܣG�,&_;tt�[�pa�*�A��������`�Zj���V�lv�F=ET����5�����3z�ɘ��6�QWG�g'�����ҷEDt�u^04<i�N�+����̇�3�@�<��C��>���)�������|w����k�O�ɩ��`����J���̔���������>����hhh��(,(����yg~��N
>�n@r!�$�+6����H����@�������I��Bx���NL|�������E|��	cf ���M3?��j��$�����3Z[�`;���u��i���� G���`C� &_P`�)��6>B�*�wJ�&'7���gԚ�/?������W��;���ObAb`�i�ͩ�qp��Ǔ���� ć���8�"��[@3�@�)?~OO���v�ɷ�˲a� �����T��ce$���UvKss;kT]�Sp=�Ydg�廾Y-����k>Y)Zxz���*#�lP�:����j;�]c�6;� ��
,�Ը�#��ʣ�f��ap�0������,x�BҶRRS��*X[u���a�D'r�
W��?)�Z��

�.k!ϟ�������GӇt�3xU��*t�o���b'D����G�
R��<oxd$XT����N<Õo�.���;��wo�a߰Y��;q}����i8�W���K��8��b�(�f׀3�zn�����Y	2~�˗/�Щ,�)� ������j�Ydef�����\�����]�ss�ATR/_�O��kyė�S�[���_I	d��qp|�7�����6gX��P�(.d�[o/p� �C�!�V^	�e��l�%|��F��L>pM����<��^�L%�����Ľ��N⒒�p��hhjj���	.���>3��K[[�wb;Y�R3�w��222Pki^q����C���^9��D�G�NQC�!%����-��w���A9@�޾}����� ��G� )\21�9 �n|��i��(5���9?��׸ #��@�� >D�s�_F��O -�{ �_**(�h�Z�kj����.3%��l���^���i�@g���@���� 5;�~��B��L�}S�������6QL�
��L�Vq `��3>:�g'�:-�����>> �ޤ�D��ׯ�/�V��y��_0bb��&$���q�ըw�B͘���d{�6��,\��{�X^��{"!'g	��	�}����k����A�,�/-ݨT������ͼ�����U7
tjf�hP���D� 2j륞�񠺉	��Waɍ�n���Kҥo��]����>3x�������k�0-d�j0\5�A����CHH�222��H�i�x�s�؝8&y�� -�c��ډ��z��v��?����SwBW�B��;��vZ���5��+++��i(�ѳj� ���rs�)�a	���4��Y|p;+����y���q�Oz�")��g�/�s���Ħ�����]�n>B���ǃ�	a�V�Cے�@�JJ�`� +n9-�Ps�"���V夣#��*�k �g

߮��5�A���o����'��$=��p��%F��4^�����pC�:W0�Sz�~>>�a<?����b<���	|:�#=\ZZ
��A�"��rrr�Ÿ��s� ��g``x`.;��v��4��W������P����Yw��ņ��'���1|8uq�E)W�I�U�R�`��T%k> ��[?��^��t˥���HIHFp��7��J�Ƶ?=�ggc{�
�!�H����������L�L���%:?�N��� ��U�JJJm�[�@��/Tj�"p�N.m3߿? d�#(=�i�*�h�<i5,
PPR��AU��9kkk���u�GQa�q�D����+����&����x0��������3��t�T����CPg�i��)Y'x��SYfx~�$����hভ��HC<�
�����T�n��P-�f���-*�W��q@
���88����~� ��֖�����~9�:gĩFD�]��Rŝ	����o@�oϰP�/�p߅xD���L�ij��ZP��om���;/f�Ӓ��{���2G��+(g�w�")혐��-I���7��d�N�Qi��9wKf�0��멩1��ȍ��}+"��R`����W�f�ڝ��R���A��G=�s����W�c��]��]��ѿ��?hR���Ōg/2��e1_���a�E'&II���SK��8�d���o��������nf����!(!!�u����H �}��H�\F5G�c���>���N"�I�y�z���r����͙����&O��-=f^_�)A��L�v��x���r����-g\�>��� k0[�"��`�H?��㊨�̓�`�m16�M(}��q��|���)�?��{0�(��G�cLN�cځ'	đFF�g����Y�R��N}:4S��LV�U�R��'ِw�K�<�~�L���Ѹ���D��h��yI|��j�p��FF�Kq�働Bb�\���$�=(�?�w�.4@`S�lu�"U4:���׀H2��mjp��@�q`h����8��f�(Tў&Z_a�{�@A��Y&���f����v��ԗ���/�pd�v�� t�[r�xo.N�Az�"dy����z����,��^���SZj�g���ϫ�D��ii� ?�?a�>����X(D<A���	Jt���# ����B�4\a������4'344�D��B�;jy�U�^N��D���L� ���\��5�C���Y��_t^�ø��~)u�vW�S�j�-8�u�_j�����H������Z�6W�H��-�S�7U�u��c�.�h���N�U�{��|����ZI�/ګ�?��ME��pꊌx��}[�����9�o��ބ̯�����)��/x�g�"�ڽ����n��R���> ��xxx�!�`b�w�GGGA9z��� �qZ8�_��w����L/șE{Ĥ�)#�T?���Q���n�!#6�;>>���W��Zʨ�^�lM���n�F��Y����� ^��AǅpY��x�P%޵kk�Cⵍ�0�z�� rmu�%䱥�|�ɭ�ly>�DU���y3F>	���Y�P�S�jm
]�)���F��O~�.�ˊ�u\F<�K	��[�k��G���7���f"H�3w��I@� ����������q�R,������CcEE��,l �o߾�d��kp�T�LV�:@d��|�މ�i{kkH�˧��ݙ�)�X��O������ stV=j@b2 |�3�D����Ql�Gׇ������~�f�
K�ۂ�`��v�zϩ�LF���-J�Ag&T<��!�Ǉ||1��R'ppp����.��mN�c:�?S�Ƽ:�b��wkKT���c�o����0�G~\g���燸�|f�i~c���1�_*(����?�W3����z���]1Y��OHhL�n�@���},���jسv����7�0�8�C��ό�2M��3�'U$=�;y۶�+��O���k6�1��]�C�G�ԩ��ld��g�s�s��zׅ#��-T!�����oM-[g�ڶ��(�ė�\]�����HhhnCBJ��K��������uyq�n������8��o7F+7U���fW��OJ�<\MH��M*;|�jF�̅�̈́���-/�;N+H�.�X�~��OU��b����p	M0�=i�+L�٧����X�b��xa��4��3����%���$&L4��y��1�B�7*�+Khtlԁ���z�4��V�꧜���#��r�w�)%������Ho�൉��q�AvT���� ��s[�+P�[V4w�x�Bv׀_�}�6A�5g�²Sߵ���;,�V��ʟe���hNNN(��5���=���𳪸��e=+��n566���_��/����r`�ؿ-n�w}����u��Eɶ��=���h���=���~=~�����=t����gS���;w�?Ў�4�)���o���э�Z:���#nn�[eh���J��f�1�cv���d�yu�9��իM�Q0�����j:::li�qw!��p�� �I�o���/�����l ��ۮ��Q�e|����5����zSS��U0�SS�,[M��_�8۹|6�A3�n31M�ܸ��biiI|!�ɿ~=�����������RZ��>��C��ڇg��\q�*�(������ȡ�p2eI����3J�����
r�Zx�3�@8~��/��`:I0�����e���NO}.�
�c5%��d6ff�ƪ��"��j��F>>'%m�x�K�3�|"" ������^� G��ag��8�m����%��z?���İ�`�:���ե��KD/6�qMg*�u	�L�.�F���z;�Y?<::�qɼ�x2��v����c@@�G����Q��L>]�t		�A��An�DDD�sveDr�iP�p�#���n��@ð^Y��mm�C��!���;-�xH����
t߯�*i{y�a�Lo�ʠ���
���ư����V[�@3�E�m��������k/�:�X�O5VTT�ȧR}�b]��P�3����u��� ��8W��0�\����n���҃0$����T���������b�i%4s����0QĹ@��T�>!ᅕ���?27g;{�A�K��2���G`VRi����;���J�n7IH�s�u� !�;%ټ��Zѱ��-!>^hpc��F+=����nV�:RL�~���P�� ;E0Z_;;Ӹ/B��ݔ� ��Lr���;R2��)��]P�l=/|^99Y��5�^f�GXXx���kpZN�ZUUUy����,v��_(�o{	��T�	���w`h�AIy�#|Z*��VU[kib����Cb�-r�x��;P��h��MdrQm�(���ڑ��#�1����#�B��5��e}�*W�P�I-//;T���� ��bԿ��h��q���CL�O�<�)�.�a5l-�J�B�#�n�f	}uef���ɓ�/_>G���׸m�^����ʽ��
��M�;l��Y �Zj�l������k�>������S'���E� �����K�#U���7.�����J�ĭ���f���P�}���-$咱�5o���w4��H��-JJ�Ǐ���23�~���t�KB�T�A���8+�Z��ұ�
��Y�K�DgEJ4�@o�_�.v|������H1x��?ʨ����Ge��вZ�`�����_ޝ���KN^[�%�}���(���U��G��C:f)L,[nb��+�q�B����9�|�|�I@"�DU]Bû� ���]�K7Q�v���m�S��2z��'ߥ������&�>��C�Ԕ���S���?���nR˿gg7�c�ҙ311}�mK�Y��
>�W�_S���ȸpp�P���_�Y��1R��ovvz⪜,4�y`YK�|�;c425e���!*;;[��wv.�R��
��o,A8g��<Ƨ��.�_�����2�^$�<N{g����nf��o���
�t,W��5���Ztrkq���;�*�\Ej7.Ɩ�y�9[��x���X�ʪ*����Fe��#{{{�ɯ�l�����~���V@*�Q"�k �aǅ�9��i\d�v`,lm�TU?&�ecc�:���)r��
̐�e@i^@��� ��"X�q��]XGO/��ӧ���E�V�ׯ_y,+\vۻ_0/#���'��zwczc��!>�N
�:�cr�W�^���d�����?|�@�z���2�QAmR���KAv����i�Jp�u]==�eB��Klu�����;ٽQ�Z@gv���%8u�99J��7i~�S�� �>�cVW�}<mԧ�����p�(w1�����������v ���A����<���GeD�300���
�JI�+(�F�����]�< XR��x^�$s22�f�������8چ�?������>^�_5��O,����:���/��q�;a�s����'%հ^3��M��^/���B�p~��1<<\�0C ��գ�Cp���MB��]��vx���e�(�*&�O@`��̀���({��z�Ӌd���tg{�����R܇��t���췘���۹Lu9�_�K�׭Ԭ�tf҉dn��#Fk��7,�@��=]�Tӵ(p�+�>ڽ �г{G�(��ל�����ڦk�Z �as�2���\>�F�揁_���"����T'���`�}��wgq��|xd� �)���H���
���V���辕���c�^^]K��)�ne��y���� o򪘙��(q>o�9�֦�����I됒�e�@�y�]��3,:#�����_!EΞ����n��G���h�a����w����X����H��W��	\��������qom{yh�r~~�t5(#H��z�0�=�['��*KJ����ކ���J�R�@ ��f���➻���ڞ�'�I�4��Jq��K�*L�k�]���3�����!!z*7�V8�t@ 1 \�a-5[�}��49���� �GX��x�<v!B'� ��m����O��bbN��;�Z��%'}�`�����l ��6��O��ݩe�i��Ģ��{g����ح1���)�cb�e9��vw]Χ(ݽ�/e6�u����Z��"'5P���E+�jb�3i��w_/*+z�)���T���qwu��V)@z���1���1��M�&]�0iag�T��[P[�}	��k����$�(��缼���qK��C��G7�q�
1���3 R����-�>4,��x�����x�����	�����f�9
	�A��[9�>��RNá:%�].��M�=��ƺЋ/��4K��_��Ȃ��J��110�%ຖSo��?vnDeꚚ�36@��m>B#Ζ�-o@�w89SS��<��}��Pl�Nd�Jϫ�`��ю�)�J�yî�yՏ�[��^�����9��q���:48�K���Ӄ���(s�sVZ4Ď��*ć��t��ڑ��+�����-�>2=�_���%�6F���3x���\�wV�#��R]�q!V
���]}}�^��qb��
�[7CBCm{�����p��AEW�ͱz�\����n ���98���#1g`�����������	�U�"�u���G��%5=&����!/�����+b4�7mk��E"ٞ�@�V��^���R����N�2�����О��}��Ǿ�-�9�x.\������}�疱����������+Ҕ�놻���gȹS�O��k�I���C(������'v��!ِ�po			U��[���z�������]�C�Lʤw���h6`��/���%�Ź� \E�nh�
}���p�|򮶌��w�O �yy@Z���v?|���Z��7���/ ?溣�I���?���+k�j]�����,���!3�`Z�M��mh�"���~�ނ�y६�����p]��R���Խ��e��K��W�����X��G�G�[e]���_��"���<=�(�D�WO�uq888� ��<�Hs�� ҷ%9!a9��7vpP!�����,4���ի��:I����ў�^�;P��������n�]i�I�mEF�當ѴF�x�S�������Jxe��פl�g�����>�	I*?�j���JO��"J2���Y_r�_:��MW~{�"þs��Om����xw�T��E�G�_&8����v�d�ͧ�Adp$v�a�����EiF+��������q��p��JKM�	
l��'ǖ;���AP�=�*�ԃό��-C5rDK��k��z�r�`�1*j��q�Og)+��o�����)=Ӎ��4�zYR>��I���x�b�bP�5���`�v�L�P��7��'yۉ>�v�=�(��ƴ�������K�4��4�C���n��+ڶ���ͥ��'���V7�J�w�wŻN�rZH,Y�:��W���3'��*����Ƹ��<<���CSv�gS�
����P�`���J���������;{������������;w��2�	�Ql���ж!��P֏��4BB�>��I'�����^梩����+��*�w7u����<�X��{֕���@��}�(:��ܯBz�MC��a�d�P���݅>:]I��V�]'��:o,������NHG�6R�R�wqM�]��oL���)�����ڠ�?߭�޵OG���c��Q�R9HC���HP�|�(�����a6�6��w8Л�ח�2��^����؟ֲ�+�ր2�t�M�D$Y�˕�U�59FR��P<:<< ��$33�2�\�j֦�g´�6��F��g�%v��,�Wv�y��.U�،{ߙi���]���R?��h�;\��zܧ�eu趪�i�2�	����Fd4h�$�)0�E6=�ĥnى�ze4�0����k��Ǆ�����q�����HϬ�	�k;�cY��g�M?�oE%�M;ngGjY�~��ЯibUѽ�+�?j�ۄ�}����Ɖ�o,�/Q�F>�U������՛���g���Vq)��n���Yn�=�A�)[Z��O0��a'�����z�a�S6%��SS�Z��\g�ޘ���ld������MG���Qd��+���}���`���6��@ɼy���
�d�]�>�!���^�\ueL9�pǤ�PQ�q�L��Z�O��^���CR`P��dQ V�)��v(K���|a�=�]cWHWݫaR��k^����m�p���'F������1,Ck�uڢ!K���ʒ[\G^�8�
���OI�fh辙X���ۣ���)=��A�R%�L���`�{�����V- o��w���6Q�hVN��6hi���W�Ū���3>�5[�x���z��D�\:�%!$H�&��E�U�1�7�⊈��ŢW<�de��ﭶ5�zxR�m�M��ɧ�鋐�Q�I��a<&%��aM�2:�z�[V?�_�1{�i5z��W���'g~}��z˧�j-Fi�#��o���%��]���1�D�긷^TT��`tO�U�/>�>�kR�4"�n6"��m��!/��-\\�r�[�*WԒ�S(�'.[���4Q���p��fj��WH�H!-�z�<������{��
��p����]�*���G���� 2!�K�?���t�r��I��_[��u��`�q&���9Z�e}����k��W$+J�v��'�dKc/N�v���#N� �!͹�dht�z�a�l\\\-(�m����*��Jo��9�ܹ���9�p��7�RTBF�H@�I������x-e�����_�qչ:'?'u&���b�W�e�1;v�r�j�!�K-�=�W\z���]��`�'	v����E��qlw8{�a@R~�ք��f�����U��o���K�K����X����]K���q�yRdw��@�r��$��b'׍:\_�%��:��y�BJ�fSʤ�i�9L����r�
VTtw��]xD�ށ�Nn�Lt"������!;���pK�&Ro�>�d�{=~��&�HFFF����W���~�-���](�������7o���ꮆ��C�O�4Ɵ�K�[�N>x�	�1j`+i�ӆñ_�0Z��-��ߊ��d%{�w\�D��li�D|������c�H������nu�HE��p�� �֫�F����R?鄶6]I���J[{_r9���a4{���XP:&)����۷�: �����A��t�Rv��<yR���Р����'������Y�%��������g%H�d���G��;�z�`{�y�q�g{���4��h�K��/��>##V+7�h���')n��������QFZ8�k��Z�(G&�����q,��x��Cy���|���_2�0!H� G�r������d��g�+��F�s�ӭ���b	�<9���9P+��*/9���|�`���߿�h=�2Ү��i�����T�!È�^(�{\ݞ�^�;;7�ny9�{v�5�)$"� %:�&55~� xx���/5>PL�V&�6Y��Ew-7�Z*dk�v�[y����9� ���9O<+��|��kV��#�|���Y����=�׿yX&0��H�"� x�X�Nd��M+ߐۭA���l:9�0��m�2<��Np���m��E�tE��?�8j�x�.��Q�|lc���
<�W��zn	���͝�{6v����l��F�1Z��(�3Ő
�qG`}�Ny1�X���$'';ΩN�X��ږ�,�D������O=�-�FF�q�:�m{�+�v���YцN*ͮ e�o�M��]}�S���P����2��Zl���9>		Q���-�9{�!ہ����AT(�v�pE�)����b����< �&����7�a/�BJ���w��������u�%t���
^&𛿮o߼:��x&%��L�Ig��Fq:����P�[)EB:D��c)�D�������s�\:޻�w�e�Ýy��y�3�-�j@�:
Y/��c�jX>����nV�!��(�t���=,l�g)�������W���+4^��ǋ�b��wg����Yq������^'zID?��a�L�����S���
 h�!�����-�y�EՀDZ�ϐ���Yr���r��"uQ���J�4�V����y�kUe�uyF��!oG�.�� ��hUA��vvvVfe�j4D���v�M�El)���;�h���߿�?�̑r�
A;�i,I|��P�
����C[��Wj��TrQP��[�������X�	y��:8���1Sg�6H�-�SW	��Ky%�7��Z0������H'���2T�̊���?@n{��u�Ħ��E�r��n�Hv.�q���rtLqL��+���ps��*�	��C�Q%BJ� ��
���e+Fs@��
��$4��**fb2���cg�<��*���V��=BnC37������;v*@����-ݵ���WlTڟ0q�(�mY�Ƅ��*�b<��c�+��o�m)��m��H�^�0������f
 %Vx�^Z������^��N�G�D�R����D��kg,%�����/��̟���>4m��nKQ�K���+�� ���t�z�ߣ	����5��������!���w)�YmNףt�pKC�m���T/����%��6L��M�EO�8���"��]��-�ւ�N|��b-�6�x6�z�����pn�D#�@|���9*���+�h��_(F����Y}��W	ˤ���A��jj��z�i\#�8��ꡝ6�Qxm��x����9K��1P�r�����BG'nM��e����4U�)��W������Y�����?�9���|�	f�ulb��h������I�����(�^J�����}���U�����8a�Jsg��[!H)?,�ˠ�R ���
׳�w����Cwҗ�6|�Q�{Z�H���[;�$367�T�ń@	�-��),tS�g����o.; 0�%��Fa�θ�?i ���������\�݊.��w$����<R7%�jH� ���$�i�5n��&������1�!f���L4���bx�V-0������{6u 8o��Y�dBʦu�0��\�����#/���w``�ݖP��ζ�#�m��x�<�9E���c�xK�����9v4�>�sk3��=8<��VH��	����A$nk���b�6�d+���~C���{_M����f3ZS2�<���>��[4��V�*�Wv�i� �u	颦��A�=��)?ö,)�'Yl���߃�	���� 6M�}����ų]�����!NNN	�:�=y'GG�e�������V#	�-�_�UT.�BI�u�<o�Qօc��
**N?��Z�I�ذ@���-\��X,�-a��l�%�c}-��fǲ*�eYL����_�y�>q�<�Z��������4p���ѻq�!����b4^�v��iڊ`-Op|Bu�t.	��t�e�T;���RR��^P����������3E�����|h������(((ސA ��`���$�RVR�Zf���	XWR�l�E8����4�5�=SZ�kae�*)��N���$�{���8�NX��S]�S[k�e�ø,;�tB�L��$�<���ԟuJc�!�/�U�A#���?4�웕�th��'�خ4���Y��g��N,�^	�ۣ����}�{�%$�`+�0g�Ȯ�ؾ:''gzbb"�bw��};Rڴ���� z+9@X#�Zow�����	l�^z��Y̖L������Y(�!�_�`���泭~��ֹ���|�Z���^5p�( �"��v��r
2"|ӻ�k����j;�;���:,��6���*��#P���S��V�\�䓜P�)!�#�V�=+�?Q����f�/тƣε&���������Y|:�(	H������r�٥���0`^�orr#����߾}c�����A}�;,�edLL����25/��Su�^�����ʥ
�Z� k~fPyTTT1����l@Qv`>��>�Y�-�_i&�9T^x88�����=�|��L��b�h�W���h�,8��/m�),v^��1"Z��hd�)�,��}HL�g��-��+���a���B���0Tv=&"="L�2�XI����|K�ZYii?[�Q����k�W!�p�שּׁ����^���������-��ׯ�ͦ=x�����g�;����
q11:�?{C�QQ
a��r��hQ���B'!q���V+M�*7hj��A<�D��Z���s��
ޅ�+��r,r��;T�|`Q���;1��4�������5���M`,�eeڀ/Zk�����<���TlX����V��I�3T!ci�7�+��ٛ�iARR}1�ްb���'l�F:�D[u��Q ɹ���49��z����AFF6�9��I���@��DEE��mq�r��T !��m�D�o�D���
�}�����\�Y�@E��D��iI�m9�!�1��ڮ�{s�0��J�Zq^�����IV,���P�ݮ,Ƿ%G��oV��WHT�N3�NP1�w�����B"9�~�5n��%� ���O�~��=�]#HMmU�vP}��Q~���S��srq��A�"B ���5�� ӭS�g�l�7��*��[.$�4l��T��^y�U�����E���o|�����kä�x���E�\�Ssr�<�p[{A�?6y���tU�pUm{HC����_����S������z94�U	drg;D0��uR�A'j:��͉������
�~^e�������E;;;�H~)��S���Zݏ��ﺻ��Z�k����N����@;;;�悂��`B��zn�~�h�"��D���w�>K�5ޏ�댠0b�Xz�e�Ӎ�(+�����6�=OR��@6Cw�U5����WC��30�,���l�ۅY�"P.���EX|z���"�Y�`6�î,����p������zu@�n"��Bۦ��>�	<J#�]]^b��U�)(�~t�a�B��YWD�ı�11�%���HH10��B�n;+=���K��6����l��y2J���[I�PR���y�t�מ��MF'nXI�9y~@?!"��Xx�K�X��!����M���$������c:��a5�PҡZ�;�ߑ�f�F(k��(1��6�5���"�&mzz:ewwW�~�yi[��<��4�p{�P:��鑸Vw�)+����Jh�,��l�u�)���1pp`hD�Ô�<�D��Ѭ2(��JW^L7<�#��(�z4]�w�>B���M�N���Lvد��ei����*���`�; `����U�~����p�bv^.N��~�֬]s�p��b���S�*�{���Ӌ$W���e���|4�k's�3�NCl���`,�9� ��p�4��Ĳ��bc�v���,  ��C�����_�p�&HPci-s�"$_n�₂}m�5������0$$1MM�/G؀Ĩ��@���
�H�l��9/�O z��69�a=o���%�\��(�)(8C���#�y}��*�&�n㞗a����b�ݽx�.�l�%';&�������ęҴ�Tu)�v��g�������� �X��qC{{{%@f��+����#�G	5!%"��ܑ�,y����3N;�v��n+Z����֜�ڢ"U��۠�� �655]P��� �s{\�����J��#p�[az��G���m�ॷ"W�*8�BHXp�g]��,<�i����l~�5�����v&�����8�:5�VO9ۨU�Z��!��̼�s�^#Y ���X��:��LB�ֳ?$GZ̉Xې07l�&��b�� �=S�%i�q�6=�Ƅ��g���$?��z�̢�I}����ު**���XD���[���̞*��T�tJnN �=���o%�N��R]af�[��̴4�Vجv���7�/ ��IJIͮx]���� ���[�d���z��)88q��j$����~���J!�;�$��u����z�1Q���AjJ~�����R,w����6�_K�*�CI
k���U<���qüqp�`��{r�wSc,}#I�[k� ��!i��w�����.�����O��n���tF��hc��2B���j������]��q���M���^���&T^��n9�mA����f6�	6��wT�����G�|#鮉�Ў��O����8��g'�3��\-������A��&6�U�[�5�mzZ�(尣9����`��>��Q��l�W8��5�g���N���mDMm��T�\W�u\mU�X� ��;,z ��M���sg0��!��<*>��UVV���Y���&��f�e%G瞦�5C�Y99e�?�(�����Qr�Y)�/�Խ=SFSӞ��O j�����MOOf?�;���미����k7��N���D��yb���X&��п�L������}w{Qk:��Vu�v%�Hi�'L<���o���Nz&��m'��2�#��'��8��f@PI�3]Y���k��{�ڣ�{Ջ>��h���ʿ/�3�(F&=�l3��TsO�^��J�*礥U1�z� O�8�[v�<V��z>;u� 3�l�*���a?�3����U|O)iiآE�A����~b:�<�ŉ�����d�5��M����x$��yVӤ5)=�4|zZ��S��g\����˪Z����{ICCCHL�?�0�^�qF��kҪ�RQqT��Xe---����\0���+�'1q/�.i�
�mF����=��o�e23G@k�'�`B*k��S�����U'�f繚¢<P���DNq�M3r*V�,taptq+�����AA��!�Y�VPi?�C'���nA�Q�΂�+i�wF�g���6c��:x~ p.X	XR`$��	�hB+��dIa�X3K��b᮹��c�1�|��4�5VL�*���x�_����qX��ȳ��	2��gϘ>R�����[�/UL�b^�N$��S[?������-z�:%{����y�Э�%��1q�}G!�qExP���#
�_�@U��r����)*~Q��z��sE���&"��lH�����T�(,,dƂ�e�fb�o{��!LD�,R=OE��hZZ�b�4�VN���U�~���{�*F۴w�v�#ɤ�44�?��LCx���3�3���:��U�F�L�V��=�U9��^jl�C���P~�?�[*�mN�O``?��f�G�� eZ�iK�˃�[	Un�+�|+b�ŖRE��:m��'^u �`��]���TC@�� 4�\V��:7�4S
�~���?ʟ��Ϋ� �����>���H_�l+��T�Օ��NT�o��1�f�M��㥤
�/#5פ��߳�*Nasy�~����\PPY��-�eZ���aXk�h:���o�� �8z�����~�����B�5���#��شj.�O�_�j�<٦���й2l~�3";`��22!�
i%b�ii�����ͦY
�zm���\ে1����˛�7�ۼ���+��4HP�@(Ժ2��[(�=�N ���,�fH{��88l���g= ��??������������� p����BkH9��WA�S{{��v��������{�����]L���ߤb�~ uU���#Lj��/^".�\�%�*��8k*�����p�h�OM�g(��Z'[?���trG&�uz� ������-H�GF� )�E�����J� $$%��r���-^��r��Z��\��B�P�� �e�����k�bY�bS#e�D���|�qZr�C^�����	u��iP��Y�L�3w��+�#��Ʀ
��ru�Ԧ�ȗ��w�a�?3��4�"�}��]i�fK�� ���40����zj1�k�Y.���}13;@�����!q���V�~7���m����^9|�b�t�:$EsssyC��4�P/���1�n wU���^���71����Yde%���~-Oi���7�ѓN����e����Op뛿1�hhOHA�X���ߛ*-�:�Y�����ܧ����m�>�yZ�+�7z瘘��t���7��1�Jޟ�G{��R��y�I)e����w����S]���\cɉȹ�����^�f�b���ԑź�^ܞ�nU��1+�cg�۲�$��i��)��[�Vf��6AZ$�7��<�֤sG*߀�EG�*��Rr�_���_&{�:O�@ļ���1U3�Z�X�_����2��~���k``�~��hp@���@ �/���U���-�~4�:^� �|g{[V����h�G�����FÖ��j�&����j��	v��+u�|�?y.���(��o��iIi��٤L��5u�| ��m�0���}(6�~y���sei��O��P�R�/�/7'�1����c�zK��<�ٹ��0�;�T��vq�����J�QR����=�.�	a4�w����͡�HB����{��☙�&&`��y	��Ѫ~}�ꃫA�C?�ٙ1��ӧa��R����-��{^2�f��!��Z��>LB�]e��f{Q�67=A���@�T�jZ2�ی��_��c۔��b�l��V��ů-c���>�v�f��>�]_/���(oU�M�9sF��*;;�j��W}�N�9������u�	����DhމU?>����ԾV���
7O�t�H33E &l���qBI��z�w����v���_��w��~�j���Cj�- d3���`�֥"SD����Y�O��yq�F^<Z�'�����	F=z��_DA""�ݒ�h@ڎ�z�ҬԿ/�kr�薒�O܍�ss"Ot�Fo*sJ$��Pw�42_\�^��q�z��{������`X��V;:\����y�Q���gS{�z�q�v�����o�X~��w�����5g6��q�N��'��̀���Qq,R�AH�Ϣ�><�%���nFN��/K���v��#�����eCW�|�B#��,�����t��PB���j�neoXGB-�x>!!��r1x��(e�Wx�TV��yNl�"/h۴�)�nK�gBP���>�%����Ͽ�T���`��V�sˁ$_)m00�������7,��ڮ�m! ���P)���vq�0P��<��}xN���(,�3�n�Z�3�n���&f�R6�V�}�V����������a��;4��qgF%׬P�4|�zÚ/�%)J��,�Y�Ӏ3"3?���}]��H�.Փ�'O1����D	[�z�=.����[�}+���r��~9n3�S��at���y�^��3ePP/��v�F^/���l�C�� m�����޼����}��˔��ܰy�=�R�1�즸2U/��A5�~�H�r�$���~,UFEE�������Ӷ=i��]Y^�\��b]'bafN�][{��5�(���L������߈A g�k��Ikŗ�'��.Ǯ��L���ʴ��B}�Kjj�ut��?rr��ˆZ����AFa����]yϛ�`�Ir�A�����o`nu��^�DҒ<!�J˄��ƶHQV��Q���&
[f�+�rveN��3]R^��=t����,���Ub9k��Z62R��@��e��9�{Ƭ�~�8�<u�{)V.�o�w�����0��j�C]w��Ϣj?H��c!�+���\�ƽw
��a�7�������u훛H�'�EEyr��o��ϖ��U�\b��	�K݁�|Z�U�mC@�㶘}��(EFF�e�ؿ}q[$##U���B����T���ssrNjBj|﯏�xW�E�|[�3ssK4�m��(7���c�\���ͯU2�`�}-�z�����<B�e�ݾ���?#��c�w��1OG�x�r�Ck�0(�~��9��d.�<�]uMl�[�ce����5���_��T[/��K��e����rx.��!E@�I\+?�	7���7=�~!d��XU���eNG� <5�ύa����!��������p@3�i��BO�ʃw?67}&��Dec��کc�!EN��fh�f/V��ҧ�׼��[������D_�������),;��7K~�7�jjbT���.��0E�M�"����P�k�F� ~Z;<�~��A?�Q�.��bq��ť�8o!�}	��xzz����G��*f��A���[~Oǒ*[Y١��>�"������U����T�R�J?]>}l�w7�9��Y�+��HTUU�f�Y��� ��Y(��S��,PbO'g���BiAg�ԳVJS�����,_�p���$�ڍڽ�����.�k]���;�j���hÚo����^��r����x�m� K��dI�,�.K5T�<��}�!��[�f���~�+#��e�Z���m�y�`mi8^��Z�f<|�V�2����&�����ȝY�{�%5-z��.����1��="�U������L�;�l�P���:�/�}�G�$tym����-�u�'�ru_vaaaQ���Q����s#D����w9��f����_%$�i��������.���_��"A��)x,�;:� ���#"222:%��;��y*�����x+��h����V;��bAaa%2�L����۹5�A������)�n����5�y A�Zp�D�*��r"���Ly4NLkm�~�h.uws
���/��4~����:���|E)� ��\�E�` ~昌���S���9J4���~���%Aɹ~����f|jHvqؐq�%>�Ht97g�c���J��!�rK�'	

�&`���7����3���ޟjeww*����~�D��A��r��rэZԆ?T٤���]o6_C�5ȧ�)�����zooI-�I]zt%�l���?[Q�ޘ��]�-�`e�O-6�ŭA��������qZ��pf��ߥ�޴�9yQ�'�D�|cc�|�G��&��B�����v&6v�{��?{JJJ�e:��X���띩0�Gn��S�X����.'R�����A�r����O5J���j��1��[�rw8�P<)vP�%�#��W��o��`��O�vrH��Rn�Ҳ�dM�ޮ�i��Z�B�A��j�c�u8����1*`]R�ŭ�얪T�x�c-#j����K4�J�� t(�S�JŲ$�*&(�:�-��KLO��R
�%D/�ͯ$:=[׽-����H&��{�M�f�C+h��bq�}��xŜμ�ƌ�.-��ec"��e�q`->U3:�*`Ua&v�8*�#Ε4�c#u�ٶ9p"����8�>�t�u(LsŞ��6��_�/2�x�7�y��j40�Y��&���V?��ׯn�ݿqf|��e|�G�(��Hkkkk`G�
z޼����Eti�`�Ƽ�>�V���;:X�:::�Z���M�:����O��OG� ���S�b�~;����F��}4�>Al~���	��ҽ��^���1!Mt��O��B�<��9F��OK���Gw���K�OD<<�O�{6���C��d��W�f��k��^J�笂��"��J�m�|=�oq�������'lg����ǒ�ͅ��c��8�Q�����E:-m��z.f�v��s��j!ڵ�g6q��/��3��c����3�[��*#�6S�O�?�
d|���I����I
	�<Ǧ�fieeU�Z<;��&:��m�Qe4��/zy��6{N�IDI)4�/�(�3	Y��\��2�qs�̎C��)J~�acb����Zw`jSRQ���g��)��vas����=Z͘08
�:ʾUb2MI@0��AT�-�U� U���Q�?QN�\�]o�������B�]UTZ"��̒ƄrS��n������h/-?7�9�{�h�^I[�L`�^����ԣ��tE0�x���J,M�8�߶z,/��*�D�*��������h|"}6�X����8����5��&!a�+$��`����FFH/�46���/�ߠ��Q|Ͽ7�� RW:m�u�ʤ�Ռ�n��W��K'&q� --�e��j�gff��z�I�d4�_���j{2�)��t�;P�H������E#sߔ���oz)v~~�#V��=��2b�Y\�cww��9�������#�ש/��#餛��*[���(5������XX�zv
�?%�b�u�Ə^}� K��D��6��"Ʀe�~�����9����2�-����Z�V�pq�J5X麿���[�p�z�X0�[�99�$>A�!Vg��J���9�e�=_J���r�p��>ۼ��"N�h��f
��{!��r�D��N�mN���tƛ>�D�}������%�� �������;a��V`�^w��ļ�>�����ʅ �%�O�.h5B�ll�*���ʸ�I\��\`��:;[xo4Smff֭V��Ei�<&= h__U˒K)�ͭ�OF��.�?@ɒL.���V��˔����f���t�X��\Y�������ε�3w���[
�ľ���:^�_ց������Vġ�����_ȝ.�E&������w?ѱ}\cA�2HH��Q};�U�l�C����Fp؄���}4`��h����

*Q��w�"Ad���O����+��*��rh�?L��y��+��'��r�^\���WS�����Q΂X�a~�5�l��ß��t��ˌ/�:�G�}
�j,4U��mz��O����ϧ��Ԏ�Lm�2� �MK:Z���^���^z�����֎��_�S��+�w�_��������������a���a�##�J�Q<���3�3t���2%�0!!��wQj�T���	c�w��sbE*/-�-Ƿ��/��y�A�G�5�/���Ď$/& ��WsPӼ�p��l��q�w�/v�Rr����qh�;#���ei�p�ͥ����Ke��Z��c�<h�t�`�u�@% Ќ��K<����e�eƶ��#|���?*����;��^��K6���g�,�v�8��"�����W���N��aK�	<	�]^���U��Z�\j=�r`�O��d��.Sߕ�,��	ϯpU%�r����Kv&$��k���5����?�&����|��"g���K%޷o��o�%&&��S�+�~�G�=�����߭^�R��,��GG*����t%��2�f��@%�V�	{Ⱥ�ߙ��ݏ�P�$��̵���Ch�fbb�������г'��Zb;���")�����Ә�Z���v;Z<u�� ��ĿC�X����S�{�О�Y:�DK?2���5C���=~8�+�zK��ko$�=%L(E�I���z[H��w�	U������VvKn����1�|�͡X�y����R��=0��0W���J#DL��$�d�/����~-��/~��C率>��&#��X0˥��~��dFv���C�U�bp��>ߡ���%�kZ'�7����]��ԙ��j��RR.�>Λ=���Z�ybV5	���x]�婩�Z=��R���K�M�`��d�<�ؤ�����o��WXT�������^s$&�j}��tT%���t���cf�#o����(,�ɩ)`��P��I�Uü�%K~��Zi�GI!�5��[y�g����p��J����F�V�s�X?j��p�W� ,���u�I�e�맞�7��ǔ*V���̺8�%��y��Hd�nQY����6���Ģ*����0�~�k�ac'������i�.HI�X_��nYV,�JO��xuUw3���!��d�:����F�U�iozgWn�-�&��[�8,ǁ���F�'���J����D<��(����� ͱV/x��0�c~i����
bT����y,-y�����)�1�uڽ��h�Z)?����^A��M�\��T�4yyyOOO�/܇ш>EMQ7��%"�5y��"�Nqu�h�oN�_f��P^�aq��KV����J����c��Eߛ;�@�{�7�cE|Y������nLB=�0�1��9�������<��n/��WD�݅uHhi�_�a P{���M0��T��W,�,J䲐R��8�yB�2��j��ӣ:���o�ّ��m��y�/��K�jd`t�(�Foe�1�7��t>ښ�,%P
�Z�JFIiy�sMJI��b�� *��ܘ�VN�h�xh����Αv��/T���1���Ej�XLM�訨��%��ci�rrr ��/9]V[܌#J��؅�<�`���ǣ]�>]�t��:��U)�������v�,ƾ�;��O���f
���o�
�B��ٻ��(ѐϢ �{hh�"�?|ֱ'��o�Kddd��X��kQE���?E{/������y��D)���y�E���,#$>)2����8xot`�$�Ӧ�������.������O��V<m&�#��H�6�l켯���$g0B�� �'&K�ZyZ
Mx�E,�G�W_Ĵo�o���y��I��� �ąL�_���'��P+�]٩�k���#��%�g۷�"<�����MÎR+U ��g��Y��q���� ���>H4�s�UϿ�B�ߘ%eϘ�Q�Z[X[CkT��@H�3D����J��?>13���l{0� X\���zr�HK���x��ΉH*�o󋋴||y;�� �׿��vRPT��f�G���g>�����"�`��g�XXX9/m�$$�s�D�b�GD��-������������
��HTE�
���9�zqf�W��h���e�<�
N&$������2z�{�D$ `�_0�at\Z@�֯H�)1�y�3NPEӚ���J����O�b�CqG\��x<u-3�9D�K:Ji
�^��s���a6Ơ�l���b�%�WOWn�l��Ջ�g7n�\�)/� �L���Ђ��/����Lxxx�C�V<�
�0)5��=�"�� �
���Y�l�����UB$dd�j��FFZNΨ�+�.AKF	�:z ��_��U}�К3�I�R���������T�ZJ���в'���<��o|����ӓ�rƳ&���!���j�@�8�p���/K��b��X�CU����n%��0����d�B+���C�*C����� ��:;��g��^D0�>=�HwgF�� ��{���D$�*�y���N��eC��QY Ӭ�5>sj�5l]؎E����	�.*mN���+Ő���8eВs$�	�������/��m_6��&�%��!`��#,b��c�F�u{�7m��A�Z����Y�]� �O?���r� �{�Ϟ� T;��豥���/���<#cb4G�J@'ui����իyxt$���?h~/�5TŸ����j��y
�ht�k����P�	��|"�N�Z1������m�s�pfhhm؏0d���JU�����ü\6u🄗I>4�]�N����9ե	�� 9�vC�d�p2'Bp@]KJ���U�V�����Ƴ�t2��V�����߳[�'((F��;��2lyz�;�� ��v'��*M�ҵ�q�Y�#d�*}���ۉuc�����>Ly���d�wJ�F�g	ziFqDx�?_h�.0��`q�εM]|�ܵ�ˡ�����s�룿WП6DIVv��4��Jމ�1OSK�'�A���oߊM��}r�;<4����|�]716�$�á7�xP�kt��ߎ��z@��Ꚛ�B�������\��A9�%�B����`���V���cbaYk:\�?� Ϡ��]|qqѮ��̶d"�C����_o�QTs�P�d��.Yb�K�<������q֛E���2𫞎<U��E_�nC�Ӯ��Mc_�/֕�P��u�^��{|��L崊�t��-�� H�Q��GvAZ�$w�/ަ���X�ƣ���#'3G6�V�H?U��ם�������D�~���������v|�|�L�pzw��_�QR�� �~�v�nN�*�{\D��݂��8ZnH,9����v�1̘��O�	���7�?,�$._�f�ujj�q3��c��N���̀���jTn"����i�������[��+/%�OB��fR�����#���"T�/������ "�o޼�,��`�>h-R-6��ޖ8��q���ܧ��$���BBAa�/�D�����oo��Ӡ!��%����$�w�cs�#`o�� A��9�����J��_�*��8ב�M��ſ8ԥ�\���X\8�_SVopo��}v�S�VF�z�ޚ$Я��g�ք��]��)�-������`O�ޖ_��ֺ�O�E�p��s�2X�����S�#G$U!Р$`�tN2jU��Ǧ� ������&M�w:�/����.��]~��1G�z�Hξ��?(w�x]g�T�������и��s��ۋ=���j@�ei�4�$n���kRRR�njn�;��JO���-O��Z����˪^��k�Խ��"y��g�|��|���"q3+�f�n�d��4x��8�ä�o�i��<��� ����f��rT����C��Ҡ�������P)k��&9�E��/n ������ϥ��{��G����Rۻ�]*r?9���d<.݊؍[j��~�|�	����̜3��giHT1���VOY� �X�m�kP�8�.1�9ޢ�-����ww���RY�9����l���)NIf��$̂5�"a�\�8˥��w^��v�^� �>�]�|'<r�Z��{�@(�C���V�׼�Fc&萁����یy�u��P=@ݏ7:�����@S���[�fj=5�9GD��������
3���eUg)�m���Kw�IFh��G`)����"����<Zm����6�3�V	������������������r�hB�/J�W95��x��ϳؘ��~�.K�I�J�~DZ���X�@ ��<{<q#�E;���+�^���xii��x� TBOMO��O��n�a�S��z��!*�*���K���"�d~��Bzz1[�p�!b���Z�`r��=)�Dŵ���)��HJ ��U�^�"��%"��I�PUb�
�Uo�\%�N�3^���=�JnF����]J��%	V�M64:Z��W	D�Х���N�Z�1�WvV�%� <B)">*/�	�p��\��?9�L�eq����7���~���l�'R+''���l��qe�:����j�A�ʖ~œ([����������ې��x��2a��=�\����ރ�����7
r����҄��k_�鿏������*�p:��� p瓗���#6��^�f	N�� �E1	I	11d��^�Y�H��i�/����J���rQ��GGG�E[w�p�����������|�,(��[� ��s[*���Wf�z՘��쯍�����ey��s�@��dJR/*�^��K	��C+N�t	�ce�g	�H	S��=��G����Ȧ�n���+��垴���	|s���B�i�Ȍ��ȝt^�jR�<��7�AH
*h�a���-���	|�]@�sm��M�������.��[��q�\>��4Z�%�=�������`Ro���d}q�,LI ᪢d6NA���t,��7 f�VT��薇s�z���Յ�Z�Yb��3=31Q���/�mb�G^VV�m���#��<�r�e��HNc���M��J��Pq��@����1�����SVŏ��۾��١N��*7&�������WaR�UF꬛c���qk�;c��FG���Ԇ9��X�ӍIt���i����o�}r���Dq��b���8�<�>�kk_#�������SĚHu����/���6��F�.`n��%�@5�Y'4=~%EO[�aM0�� y��^��	�l���k����a%��p�ҷ��%���l]6pa��{^��M��Te!�\�Gzo�O��@�n��U�?tn�bBrF!Y��+4x.�fw���	g����-���=�s�_$쪍)@DD���/�>< �"�gM�%''�s�h��,�&Lߥ	{8��X��eMDLz�<r7�v�(P����_dtw>��YS�����B�*:���=::ʎC΅�Z�^�y���>��^�����R�����T�K2B���UK���p�{�vz�=��7Nn��B6�Z�c܈�TUp��Z��k����w��O����'��x
C���-q�gA2�zCE��?�C���[�4x�����;>0�21��_��������\���[y�bS 	EhƼ>>؋>x�l�ps^4��1n��TM׊;�X�if���kH:+����)Z0���� ؋2�����iF�W,XB�l�����2����C���c��s�{^^�U��Kz����Q���_�sw�E*�	ɚ�̱�����p�O����i�'���ȯ�9������Kv�T0�m���hpymЩ��H���ʲ� ������CK5�nviiI��P�~�L�vzp^%6ɻ�������ܮnk��52�RK�0����;��k���?�kw"�1��`���4��{G#���������Zo��Di�n"--�>T�sݺt⡣C��� 7�k�MO���I��+YJ��Ö�zR+��X1r�����Y��1���+���u����޷?8���*9�˄�oȏY���p]]��C'��m%�D�̂	���A|L��!#���
%ԁ \}�2�;;x`z�F[�Ĵ���0H�^�}U���mC��L�E�d����p��}lYq���ir&=.n]�@��YgD"��w�p�S���r�����/?to7�a^����R�# @^XX�d=�ى��$�oHӳUoA�D#����[�E�}o�CH�4R�]CK�4)]�))"� "ݠtI��]3t3p�|�{?�7�JXg�g=��>Ldyf�p�!� =�׺e�t"����z�����5r$99�s���5����݁{�P֦��d���S��һ?�� s���|�f�ݺ�~Rx3�.׋VFem^%���N����7~�[%����x`�2�w�/�����obC�_?�VԺ�S����>���D6��}i��B�[i#�:�*C!CN�>��浇7���S�� 0;5'��l�����*7S�d����W,�G�B}����bc�J�#-���R)rx	S
23i؊�͔)�9��@��?����]�St1Ͻ%�iEC��ʋ[w���w�,���'"��	EMA���QS�Dsh���ݑ��Ne�+��SH�o�X�{y���rLy&�员�.���@�.e �9��[]?���T&k�J��)O}���~�`�vI���U�ؓ����{�������o���Fj�dI��퇋e�HH4ޥ��xN|����fz5����b77o#����#U�g$������Q��P�Q^���@7MG��M����j�O��0�R����;����=�GGWٟ&�3A��H��#��PQ��,�����ߖKb�3^��E.�ьl�;~Y<��+���>�*Q��y��G�n��n���s"7P�<V��3ݩ����������*DH���ƅ��/5�5�{y�|���-��<׻��j܆T�Y�,���?�r� ����;	D��?.���N-f��yX�oW��p�\�R��91�#�}%��ȍ��_/�)��慜��;���>|L������݀�h��s�~�'���]�P	�n�!!a0g�Z��N����\Z�Q��t���͙��:�k���@7t⓾���*�������g26�N68L�'�p5E"�9�����j� ǿ|�	��֌*����7zz�S�� �7(V��
I��U�~>��r����Zm	^l���U�}�������$�ŕb"��$��Ӟ�g�M[�f�4�q��h3��'Wh��r�d�#s���c`q�u���w�~��!��E��w��?Y���AD%��ށk�8	����CHD������0nI��̪�j""Fw7ǥf Z�@��͊��(<@:ˑ"IR`�:`I��2yq<R��ɽ��"�!'W�p��ҩR:�n��"=ϰ��kv嬣�ҽT������{����꿻�*�섵����Դt.�܁�x)m��H���^lnZ��[����Y��nr	�^�r�`ǵ��s�?���Y)\sc��KH�v�
��J�T�"�xG��i���z�Y�mi����͸���$  +���:v X>n��a��*�z�4�󞆍h��:��X@lyx!n�+�1]���Ҕ�?Gt���P�ޭ�������n�rB�z�����Ua�-�ޣ$�&7�J)De��R����%��H�j-�"!�K�����x�;�b��ӄ��`ma���3�����8�M~�u8����-�[��������ܦd�lބ�P�t.Gb4@ �C��,a������V�R;�^�L�������1�K�3�!M&�fS���SL4|:������a�2	T������p��9�I����HQ��\��1k~����O�^"�$���x>���	�J�2�.D*Z5��7����w){GL�77��*\J��5���ZߥɆ��(�(�(��Y�4u~���`�,��^|���&�:��\ S�aD��V������ٙ
���6�'2��z'�������ov�h7�vfDh��Zan�c���
�e��R�����K4Ow���R�|k(���܏�������'~�C��{Ҙ���q�21�d*����rz�h@8.5���#�&z���ç+P�-��~T)U��h8��:�FFzȅǧ�` �����uiUA���g{�WG؍©}! s���x��谢f.u�z�WM1P��'[o��U�a�����9���H�ﴺ<}�������.T����a���eY5�'O���q��Rس�l��ŏ�12S�'�"x�=b�u�v|&�L���ݿ�(
�a�e���OE���慑@��*�N��$I�_��xw���Z_�b �wX�R��R
c%�0U���E��Zr�k�/Q/;��+kh�}�4��G�����J�J�{��'>���ce�X�?'H1�^Qo645���`bo`�a��%t�-bMG��.��zi�����y�(8"�%qĕ25Nyxwi�V�(�̠XH�RY~י<���J�Rv�.bY|��3yB���f ��y ƽ�Ge��\��~�h	z&bϧ�3�!]��x!{+'	ۈO� ����ը[ZB"ँ��0���|ژ���W��S�Ϳ	~��� 4��@ "�}��//�z�r�o�^�EK�s���M;�W��.�mY��`�y�����7��B�����O.����&�N��rr�R������'AFK����#��8�<�|���~ã^�Ǵ��n�����Ga�H�3^r�ǋ%�ba«��2hz���򱖢��W2H�=����C7I~حa<"��qvQ��l��ծ'�ONL\���b�Ɍ��i��:ZZ�-e�,�,zTTU���ehU�I�L��m�3��{�98_c�?�����qw�*6Rމ%3�VS������]��UVUU6�%N�JƧ�F��(=��[#b�rF�q�F�=���[\��B�=yا�0��ۖ�w|@Љ�:����c��cUz���lD��ɇBUC�o��^�_ B2�UÆ'�a#�z�g9+��_��\<���3�����
��&TG�����֕ޭ�q�w}�v���ρl����}{x����,���\�D����P͒�X�������-���<�-$)I'��'?N'  ��$���ZSS�����<zQח�F�?��`��H��E�����qwwp�(�e��z��֊zűP���~�7�*�Z&�
t#�*2�%�M���=��Hh��Mt�	2�ʪ�m�<����>`RR��i� b%����@f�B�*��tf��/u��_�^_��&:9wx��[���*�2?�\��8Ӳ��`T�s���~��~KK�D�P �[O��><��5�F���ۻ>��7�j�-E7�D�������:^����Pt�	�kڣ����7��A~TkY�qy�O����÷�嚵���m��ú�I�7>J�W�>�Q޿�
z���}?�m���� ����'D�X��Q6F�Z�]L�x��,�y�hl7�^|M�D��.]���hPD:iF���l�%'<3�'α���:X���e&Q.g�a< �oh�]��V1pF���p='�Pk����Έ��BW���%Z..� ÍY��[M��m�/����A��߿y�"EU7�o�}�S8��N�qpp�'q�nlH�@��E���(8I���\��"/�����/z:,�G� Pz���y�Ķ?�֟�ȍ�U֛�����D� �*@������<�qp哧��C8N���YRZ�ǐ���oo:������3{�q�$S��1<��ϠJ-N�.��}���1QR�O�;,��R�+ƍ����I�ں1�;] 䧿h~�Lvk0e���jcSS����	I�P*wc9ٻ?Y��4S���/����QQPP�K��� �򌜜x ��h�����k�8�3�O�]�jn�Tx�FOoU�!�&gi��ڒ�����Y���G5����� ���*4U@�bB���F�!��!K��y��;��kϾ|��o��]|"���Mv�syMܓ��MVT�}PJ㏾\�=��v��u�![O �4R5ѹ���dqwYM@f���/��f6c߁�(�8�j�����A>�B��A�����~3�`2?!,I�'''��I��>p01��yJ[[�H��400 d�(��P��:�nw!�qId�������/��E�5}�d@H�0:�ڱu�p��k^�|$r���W_3���_dh}[Ip�5�\��@
�����F����s�2�$fu L�'g�"ڰ"?{)�5��7�fB�����c]K}'�)��T�Y;k!�L��y�O~m⃫��F.ߜr�V�� �^9�7�-�#���/��"�]l3Y�7/G.^6"sq����tSysk+����v=0599�`�2_&s���#�$2�5��B>��v��<xН���>z���^;0w$0��3?��jznu��T�o�UjKd6z9j	G�öx�]<"�\^���Gq9Z[��^
��S��y#��2�E�<�,��<��o�_��$z�|���W,���	�(a����T�,��|���,��^
M�@ݒ�Zy�k=��'�4�D�	��z����:)��nG'���z<���a����CMmf�Uu}�а���;�M<G^m�c��j j�SoO4����z ���Im�K�Y����-�eZA??���7�7����C�K(�2���;�vO݈i}x%����e�����71�e�SMӌ�GytK�oǍ�
 n}YNwz��V�]�Ʀ=��`}{˷3c�y�����-� ��%#���1�Į���C��;L�VU�p�L�����F]<ɓ����!d;����%֡uV�=��3���f����<w�))*��u�ԕ����7O��9��ٛ���]6#H=(����(݊p�^�?ga���7�KO��k|} e�Lҧ�.2x��ƥ�M�N��a��@�[=43$����LE�a˚�M��3�F����N�D%���	��.������%L�0��B'����)��-�����O��:$������@�,^��������0�Jj)����LFw7��\s	ȼ,�Ͱ'�d����\O5�}oG L
8���ˬ���۷O��^�g�M�eb�;��Y���?����T�ߥ���K)K�h)�$ѳF>z��z7�fl&�0�=��בּ��y��!y����]�n\�~�h�]��fq�U[<����\qN�$�Q��V������ktb˶	:�9�2=�v�����{z*�b��	�*~�R�&G�@~�9S�@F*\��(�:[�ZTh3"#&]G��k�h{Gء�>3�Ϙ?=�_dg����-kn�r}���DG�F&=�ϑ�!����I+?�&Y��\(���\]�r|y�����+�`���r�h��ǏA �G�~es�yE*��j�{�ǯ ������	�M�HpI3Mj{ox7S�2XG�v����6�ywq����mO[gB�7?]v�?�ň����w5�x�u�;>2B~��n�^�uZo��o�p�-F�+d k�r(�o(�+�O#���s�~`�{,�٨�Q5mqhg�������3���V�hpDy��h�`����&<8ޱЭ���-�h�V�[��\�|	{�������2�R�T$I`#3E\��z��ڡ��}7��h�+ЯwP�Re����$*ms�Yp�k�[�U|���6��0��Oi�jHg�]��>�z��n�`�4̤�"�r���b$ftsO���>����lKF�y��ځc�xW4�ﰥ��M�����?n����Uk��D�A4ކ|���P�糘S�X�0=<��/_#WDs
���h�l�1�����Q�>N]t0&t��s
���L?M�w�������Q�LX�}��Ћ��H^�̮�Ow�L���Ƕ�,v�km�IH{>ω�i)V��-���� �ᄇ�PЏ/�a���d�� �l� ~�::�Ư�/�[���C�̏�(�Љ�k�-|��4��~�I;��5KX�]���g�R;���@�
\j���K�s��/RA W�>�N/7�~�����iW땅Ƕ�zے�"" ����$�Ą���axԝ++�&&&9o�vߴ��ݠ|x���.���������J�W�]==����\�R'R� ��e}�D��(.��l�k_yI�j��A��i#Gē+k�/��N�l��A�����7�/ŚV�ry�`}���d�Dl��])��ڥƶT���~P�C��]�?�F�PNg��sM�fbߨ���
��$><$�oQBPXȗ�Mʯ�_�Ʒ|_��E<姿���:81��Mo�Γ'�Y��TT�j�,��ng�j�==��j�1J"�YO��?��Ӑ��ļ=����"�A����{Á��9�q o�����}K�Ͻ�Ga���4��c�|�M�9��Z�ߤf�X7M�1
��r"��-����_��%�Z�:��,�Q��~�F��$��ӆ궿�+�8��7�߲�i�PF�1�8�3GDl�y&����{X�g��A��
���i�)�S̛,�B�þ?U���:��������[iF[_��L����[�NK��m�a
&0���Hn�:8�>>vb;vp��� ���1or�g����w��ßH���0��J�@��+����?+��y�(�Ul�F
t�]o�K���E
�>�#9=��4����Ms�D����s{�;����`z���,���o�2�N3+^�(Wv�Uǂ	�C���	2��]�������@����A�LĽ�~����3 �roռ���++�b]O$	��V�
��Ս40#`r���v�)�?sbm�X�}93��Z�֢Cu|u�e���g��CF6����8B�Ab��*�4�!��VI�z�G�q�$>4��3���5����6�ϝ��4$����c\ǐU�%@�H{�ilp���p�!r��7h+c>�]"���!���{����ܚ �������z�����2Gi�~W<��z|T���.O�0���4�J#�v���?�Z����Xv��Ѳ:���pC�G!��I���T�w�һEEE��U����vF�88p!��x�a�Ϫ����{:i**j5�tvʲ�q5�XYմp�Qj!� �cP(��@�"�`{O및���1������_��R��N l�<����[^�� ���@������8�m��2'�~� >_�ң;�?F0���c7�җ�J�uv������UR��hRhD	��j�R������ڨVCf�Sq�"#T�;�9�@g��M��צ��>a&d��a|�3>>-gm]���>�;���JTrZ���k�eռ�@1-���aȇ?����x�d�TO.�]�9�-�7�Zȁ����a)x�e�.А�F��W���<;��/9q�S�+�W*���ڱS_Q1������O��x/�8��m^N)�&��V^�X��-���o����/�z<�h���.��B�_(_˻�F��O��R�#@��;숪�&.�ϴ�.�L�4���u�;��/��^�x���05��v.�bI��N~��%�t+������ѶT���sc`�x�H��Jc{7�����ź�����ղ8+"b�� �c�@�aє����r1�&Jαg]�����o:�P"���q��s��4��ӵ��: ����!��h��.^��N�@΋�:a�aP�o�&����;3#iOf:��3�2V�4�uo"��>�du�1
���V����ED.�V�'Xt7�d�.Ί׷�!TQӞ�h	���Hk�?���/��/.0�p�`��gM�[�j6�|�aVur�邿*�=p4��kԓ:�d""Ð��u�E����6�o��O�g��E�<d�9������'j��+��D�j���t�M�sM���+`�����0�$`�e�:�HuP�l-�wq��f�_�-C�}�M�n_[�����~19�1,j���Sp{,��O���[u�S��!G�hVtL�����%Lg��}P77G.�Ȩ��y��&�pB��Z[bV��v L�Y_���R埅�oӲ�`%|�ٱ���'��������!����2�$�����wW_���T`�W�{Q�:9`�S;۞�/���pQ���AmM�Y;�/.��}��9#.�O�h"l�d���ڀ-�9���%��;ͳ��>��?�%Y���sŋ6P�d�1\����S&j�@���wIt={�uh�u!N�HK>�x��A����K7L"-�	�OȻ%`&"�YF��)U�����Lp�D|VV2�`#}�$���
*}�G�I�L��3�����%%�DTL�V��H�	ђq��W�r���P�ِ:B��heC�-����hV����!:E#.|��&���T���9UR��3��AH�
�퉏F�~W/1�9d���ߢYX����U1w�*�[e�Db�����Z�(���Y�H�B��G��B�!��M",\�d8�����5��D���͞�MID���۷k�v�Ԥ���z�FG���R�M$�]U���w���c��!DAAq���1���[�Ԕ���\Y��V��{2?�� Ą��3�-"pr��ղ���V�z|bb1�N%��Rk�������׳�q*�@ͣ<}�_d���d�w����zf���l(�3�/:�qɷ�/��[Z>�s�|R�����A�v4�̮x�6�ly�O��q�d�����`O��P��xNs/Q��a*s�%+�vGd�B����
�H���.iyC��0�y�k{{��5.��Wi���\[[*ծHS��(����}C]I)�_}Q����~�R���M�>�uM1?��hDDDS Z�H6ҸL9�����<�&�vq�&wh��0�L[�SH��ʋ���T¡h��չ��o,NN P��q)�V�U&i|�9���]�S���au����9%}�_�۱�\��'Ov���� (��ɟI�@��X�G=@>d��9�|<7��;�4̪9p�s�M{����(k��r��n�Ҹ���g��ww�4������@��})������W���)x���^^�)�����\�s��/H��j��T�E��� �X
R���fdNo��]V��ޠ��R:�/���zحj[����W����p���+Ӧ���h������1טi���v.e�MLO�R�p��)Z�3��,�1r�|�j�X�Ή7g�q���93�
�wG	��@D�9�]^ް<[��x���$Fc��͠�2F6�;�)�P�	4d��'�����M���
U`nV���"	�5��Uy(���^"'�YY�m�Cv,�]듟�_x�b>-�r��n�.-.��1]��5���67���f�fA��2��R���� 0�@q�f:(��Z�D�p�԰�#eNaҜ��[;쫋w	*�yf���7陀_M9W����F���v�p�ȿ��	!U�0#�/�~n��iP4	����#Ox��X��>y�����b�����M�/`�w����*2����b��v��j0t0Xd��=�����/��������A�����G/5:�=�do_0�w��?(:���7�����܂x��M��Y�R��:�JЄk�!Ԕ��WR72:SPP�L>`r��G?Wh�x�ۜ�ʋ*_9���;,3'�q��ط�8`8s@���Q?|���#����9�X�Inp`)�����"ߘ.G��:�!2�r�P�jJ���,��.��%���Wi��݄��^˞�wM�D�����2����Gv��Vg�(A���q�_~�����j�}�:n�V���I~$��j�]��~Ә\�j}�:�7zPN�0\>�"�/�q����d���Tu�@u�踦f{�k��t�Ӻ0۟�m�]�������#�7��|����i�4|�m�:^����ʖo�sf��t���\˥�~�� �7�M�r;�����6�zn��|���a�п4�%i�_5U��l5K�te��J��+��*\:��~}�k������*��~��5#U��2��h��v:��ϟ�RF����g,���weR߱���'(�1��/B0��h�OM�o����o}((aZͬ��\��<0N��z`�h*4Q'���K��� �hW��.�6E��f��)�by��F�.�I9�%�Z-Z��K�	$�Uյ:��o2r|�@3�BZx>Y��Y��L����Pk
~*��tb,/�lúw���~4̿��V7���TZ�)�v��4�g�)dM<~:u�>?uE3�J����L[��պ�A�=WP��'K��	�@ �����j.�e\ie����he�J���W�K�ñ��B�˒��%��ɚ��*u��՝-��l�7�4Q �ƋZ!������l��#gw~t�EnS���������^���1��b�?��)���y��i^m�/�t�����N�J�������!���w(�ԛ��V>�,�-UN��jg�,��Dg�fX�N�X�s�?���	@��4��F{���dv�L���y|�
�b�nlQ��P}���3��-$4�y������8k�����N��7���A{:P�4�H�� #3�g�(���s�'�+�*$�e0����yݯC�T.<3�(_Y��m�QbЯGl�������^�D����iygc�|7E
6g_'-"�Z�w������  �Ll0���i��f�y[������ł���١��/'$;T��vs�Hau>����SdG$������ŖЕ-R�JE�����/+�e�nd�~{���̛4�����J�c$odS���@Ny���Zq�l#����n�@�M�+uh��#�)���%=sFM:��p@�*'�@~{=���R��I��d�=�y��9�#��$ծ�H�������:E��Q�)����K���RE�눞��`сG����IM�}`���tFu�P=Vs���"�h���>F��5���Ki}@/UT��X�=����6��M!y{^iR���S!y����GŊl�*mu�,��"n�yΎT�[���DNX��u�=[<���Dbf��b�9����N�7ʩ�6��v���=�q��4�n��>��+�x�#_9v*����;���e9�xM^�&ɱ��<f��+7.ɗ�A���%�v�9�O�lF�<�f�㞀�lg߯��Ud���_2oS*�1D	���:�u��=�f����s>Pl	�'�� �;u�p��"=ۉ��mxIffn���)���k=A�x�h�ϼ�Mٯf��Kp/����d������t��G�'�
�v�j�"0hۣ�P류�~<N�PUd�/�a�����|��E�0���Y��
��k���>?�A��X<p@�P�o<��~��;e��Q�EB��]ִ�����.�����,���Q���`%֑`�@x��)���듎~6�S��oXℐ��ȭ�6'�T_��>Gp�/�,o2!_x�q��+ֺ�<���7������^�����5�>sLN�Lf��/TJ�"b������U�"�c��|9��_��N�0��O��A�
=�B_��^��4���(�,�����J��o6K��I�����	�!�Y�j��Et&�j��͂����(�Eu�G�:_w�:jbV��rWWe���8�qw�yCU�ۈ�qrM��f1X�W�q�a;w����8V������ѡ7)���������ߞ@�����&��?d�凛W,����b���ɢ��W%گ�܁b���D�ŋ���x��R����&Kw�薐�F��L� ]� }��~�KT�j\�4�@��ϻy�썕�������&z�å}�螸�w]�՘/r~��k�+��#� ��s]Į�ݴ�Ui�$
�bBD�������w@ta�+9�֟�<��tie���N��Q5 K+1k�B!�� �RY�U��ܳ���0��%f�AՑ��91��4��H�1W^�����g���G�!��R���6};��o;9C�7��h�`黇�&�(���]�D�	���f��J���Yb9Ʋ����.�3���A (��ŀ�㥑@^8���&]��"���ԁO��2��g�׼��ݻ������$�&��5;�W	e��ŝ�u��&�v�)�y��<�$������lAp(�D��S��n?#G�� `���� �چՊA�4�g	4�w��s���pd�C8���j�	���Z����/����y��j�e����CI�<��U�[�r�d�n5fCg�����8l�bs��~Y�·#
ҹ��}0����=��Llxy��Mt!�͢Qz��4�;�N6llM�Ӕ_��ɶ����
��*�
��Fn�
Z��.��wQץ��� biU�J�1���6���.�5Pτ��_�V�@I��?6���V�ǻD�e��s,�Ԫ����ڛ������ӛ����a��#�5TS�i��=����t�2�|*�#Y�?'�K'�T��)$�����kϱSanr�_�mpV���?Ӯ tA�Jpn9ֶA�GX�h��Q�A��bdw���z,F�mQ5�����$�d�,��f�K��,0.�P��@ݤ�1��T��nG
���!�3�+?�9��p�E�#\���[�^R�{����G9u�t!�E:�0�j�ڇQ���D��hdzpx�\0�b�rsb�vj�O�6��b���J������J���bR�R���p7��p}S��H	U�U�fprH�wu|��rH�+���j eVuN��W��z )64�ھ�h#]�'���`��/�j��(�����ǹ"�l��Q�F�n f��ڡ�7�4�L��T�V)�dc0 Qíˮ�(Qr(5U^3������r�m��cʬA��[2�Ȝ�L�eC�����-f7���q�k�_�~�vv���.p�Vߐ� �SdU!���GV,���pj�\�(]�l̴�����d�M�)~]P�55�����5Hy�%�v��32+bp�-�&����K�H�\

?��4��}r�2-.ϵ��{Pɀ&_NlS-]�|�>��[h����;y��E1����dΓ��5W�PTϖ������š}�HP���}v6�W�'�h@�\G+��J��*ˑ4H����w��W�󅪀;m��mi,d�w�I`,�5/�k�v�x��KZ�5C�6`���p<��a��Ye��A�ƮG�|�F?��g+j�˸��VN������	d7��,�q��z��-����N穗�ow��&���M�@i�^�o��L���$Q ��Bđ�0)��m��@ȩ;���j��?3
Ft��U[�QV����O�,�D=� �!@� I��wh/����N�����?��#�����P!B��Z��$.a�D�V���gx���uc?�ppr���i&�Y�ƗT}�lPA4�; i�������/Gy<"����	k�'� 
>̒��=���y	�n�{T��x5ր�e~3Մ��5�K���A;��Z2! vGR���0{�����s\��.Xa��R#��0�xa�����ե��W�4�;6���	�h�)P(`����/��F�O{H�Aש�L��P�苭�����pA��E��W6 2����ކx>3�ؒwk5�Y\��22��tDN�x$*�o��q
����+v<y@��nj�"�+�ӹ5@<�-f)ܒ/Xy_M4}�ٔk�Uԁ�Q"jN�F3������&�ܯl'(g٘��@�q6�+w�q�����Ń?>�_�Ö��~VBj��ܣ��tQE�������ӷ�Yf�S��������@���z?���u���).��h�[YI�о�m3����� �KI��(w��Z��J(��eF������x��ʽM�t[�w����(�Ag���H��;?��6<�ә���V�t ��كq)�����79,�.�3��ʵ柲<��0���6�?�*���On2����Q�&���>�g�0Zӽ�J�fۏ��*�}�I�7nҪ�z�NMkW�>X�P�+Kȡ����f���o�r��pa�P�cq����nb� 9MH���L:�\�	�11;��`j�d�E�v��~�1<���?^�x!���Vd�=E��s2��Җ��
*\��c�%�Jf�lf�N�w9pp�A���O	�{'���~Mޒ�������_�S��m����ac�va7ш�w��ڝ4���7��K�#��Phl�����+��GD���'ʨ�y'�sLt����*��tr��t��A�b���w��s(T�/I��פ���������/���U'9yR�^��qO$�+�?�_�RnN�����~��t;-'j���BM�l�4Qm��c#ŷ���6�}4�I���.^���z�}s��#����SwE	��x��[s�2�f�H���p`������L?|N`�,����5@N!�ݾ�IN�`|J?��g��7pO���y��:]�hگ����=@��Ё�u;�G���K!^���|�t��pw���b����t!�����W����6]Q�K��*����R
5V�M@�V����uW�+��vW��W5�^߀*1���_0-ޖ��8��V
��"�]��[$N�q���1�䌮5�%+�_�ٜ�c���➕,�>E�f����^S m�Y�> n%Q�^�h�]�Ds�T��1��q~:��<n���7&XvW�G�^��q;�0}�q��b�������7 ������u����i�gk���f�B��?��G���󻎽�zI���5��
�-�bW��S�����W_I�]6E<p�z��yθ\d��:�t0垙�i�:3n'LX��v\J1g?���$HTԧ��fIc6Ȝ,�^�R�o_�Rx߶�}T��e�Bہ�*o���ew��2�)�z<H c�������z��s������F�֭��=��o�yd��Z±�E�ܩ�&?�8���)��K�lR��68Y`+� y�v�C�_X����a�T.9}wS���=&�o��^T�KX�s��]WV|�iMkB��>8{�xI~~B�Y�!P����i�+�Mp��~�9`�X�/&����^��V5c��>L������>v���P!P���7�Ө�{4K�NR�1�xI�giٚ�|���l�'�bQ��u���[	3J��i/ak}8�6�9�FКw����"A[�@A�yj��׮>�op��x\�"�}����}lv�x-q}�^vW�|Zl��ٴ=x��f���O.���V�À�Yo��A�^V.���~Q�7VtX�t��1���sE�]j�0q	q�b���hM��1ŕ�B�W�̢���:6]�tZą���\N�$<h �	1�X��8���0��E���YVGCrN(���5�u	���$d�|"B�D�%���n�W�3*����X�P!���t���\D�Ļ�Z�� �y�T���'@�ݡ���1w�eu�E���āݞ�[�S����:��{��#d񻱡в'L����Z��f.:R�*��[�v>�:�}��������}ݚ�2�7n�ϲZ|�A V��~qS�q�f{������� ,󊃓� ����씠�kf�·�{6��
~P��NNL�x�
r�j�Ϗ���œZ@12�x��mh&�l�ڇ����=���Y0_X��9�x����!��Ӯ&�s3`��g��,�R�,�Ű�{�)+w����(�w;3���9�,q[��E:d���lC�H؞0����&�K֩yݷ����K��&��^?)�� ��� �6u9���u����p������ ;%�
�V�Ꮂn���9\�o��{�%���=�I�ݾ��%�N��|Q�+n�_��z��׳��w�sKZ�p��O$~�@Ed��� s���Pj9�+YDM���K{:V��@�{ߘC����3����L&�7!v���kkh�ρ�1�����67iaO���	<s��
(r��p�2!�ۋ��ҝ��R�iy]˝�	V!m+Ϧ}{�q&��R%(�lYZ��6:!���>z#�|dP^���0]by��u���g&q$м�-)D�.�32-�QW�2��%��/��`�=y�Nݗ�G���|7.@�*����
{CT ����!�J:̥��L���D��Z�|Oг$������?}�=�����֮�g�oH����9>N�Q�.bu�㈀f�Xi_W����A��5_#!bZ���%Q�H�i�sɴN�� *�g�έ����x�K�V�����,+�]�o��e����.@~s3+�(�ZO�>+�PO�$tŉ_�X��}f����KH��l�<ȓ6y�Ҥ�q�����m|�e�����2Ȃ�����;���cKL{a�����KG/>�d{� �=
J_�����w�����.s��gKi�ÿ}:�lٝ��I�<�,�`���,��%�k׶��]��:�%b��-��˷�`V����� PW�J�A���'��J�=�����C�?�/7��-�ӿr�����%����)�gI��=5I���](T�ݣ�Fe^�F�o�R���нnf0UJD�8�N��n�[�e���� b���n �^�]2綴޿�>~�c�?~��������g�Bf5�R�i���r�����{��I!�}�S�A������5��=��p���*�\�|�V�8Vy����3�����׬j�^I f|�lra��ք2*1�s��_��w��2y���Ӆ�=����Yx���b�CO��2�[��(p͊���������T�Ѫf�C�B�� ��WZqY�B�]6��@z-&Bw���o̸�T�8EzK����"���0�Z�_[�ŗ�?�>�&��X�5�Ot��%!�v_��A�(u82��x�=y�>2�*m��p*|آ�j��|�C�w�Z�-<P���[�x�i��vbF� ���SA�W(r�?�&}*�U��KO]��f��޿��s�jey�ᇀ��\JX���e���V��쩄D5(��L�����o�����IT���نu��P�4j~k}�$��J���;������!�7��Z��UFF��"{�̔ʖ��͵/���^�ڑu)q��;���������}����|��9�Vn����HG`����t]��g�y�Uq�Z��ѷ�=��TC9�(U���	��b��j�G�����r_L�O?6՛w&���Y��I��P�g�+����������Ѭ�/ei�0!w[138�+b~�M�����2�8j�l<�_���4�E��ƅ?�Cr����8K��P���&q�Z��P���C���C'bx���g���S��䤩�7���]�7xx���q�x��*�g���	�w���{�6����G������ O�4�}�ԍ�?:��_}��{���`�M����s���Ok�}�c�u��OK;��-���$V�ho�X�t��]�LMC�+Z���^
�oP�� @T�\N2��F�U(�>K2���)����v�Y���R*��瞯�F
��`�{_�(�A�ޜ��-��=�8��c����?�W/D妺s�1�7���̿�٢h"d�� �E0�X�D�CV�+]:�k��=�^�Χ���Ғ��BO��T�#V]�z���	�V��fz,�l��b+ͥ=�;���%6R�1o�U#�׿��I�(�2ɇA����X#�e�s�7"瘵�Y�/n�&���������h~ݛ�DX��X�h�����&�@T��66����Yr1�di�A�~��p��}����.�-=Y��}�� ��̧�g��{�T���W[��/-�Р�t>\����dWec�_Ϣ����S���/�x�����Khv�!Id��v��k�{ُk���J^�5$�D����[&|��4K>Xj�I�����$`;�����k�ͤ�%�g�sO�`hEΑ�_�v���`���.i������8׃Y��P�6U��Yǁ�P@F��<T���b+�FL�?����k{�������=��rm^Y��e[H<ld�3~�<��N)���H�E��������IW�o���g�� C�CC�瞣n��� j2m��ŭ��2���0$ D�Xa7o�*B��bo�^�E��yyS���,m�$�wL��YN��T��3_�_����Ս�y�����mL���a�g+�3��8v�D]�-�A:�/\�MQ	���Q~�&x��h.��8d��٫w���\]O��| ���e%8S5��E$0�X'�!�^�D�DF8a�b��aO�>Ґ�M;̐?1�L�A�t�v>�訵�����4ش�Ys�˻z��_<��� ��G��OMY ^y(˔]:w�����WChtT!��|\γ91|����R����M�׼[ �b�݅JYB���ӿ-t�H��b1��h*��&�^7Wqx��8�l涍��ޜrV5�����=#g��Z�R0����C�T�'�"�.9?�S�J�h���#���u2e�{:����� ���n���ӿ�(@�k�3�N�L�IUN�n���D_K�q�[Py�dp����IM@��	d�S}������}��mPV/2Z|:�����v������{�OG���JOQ��{qa��&�Fb�7�����}ܜφ婤�� ���K=���1�+��臦o�qS�(���Y��U
�lB��7�Es�� �8��r+M|�TB��|	��!�K���q�23Q<+ �,�f����Me+��!����Qx����w��	�-��ݐ��L\Qy��B&��ǗK<i�݆ޛ�&f篤F�Td����:N��\���4�o����t�ɧ8����m2>⯓�.^@o�>���j�������Z�ȵ���Y��FC�����&�̑���WM��.Q��;(mR(:�è�x�t	�������S������Au��gjU ,8��&��6�r9����~���u��蚎���3=�~<Н�򚋧� Q���u���8����x��CѼX��7����P��9�>�Q��6:/�8^ߟ,3d���"EP:i�D���S�20^����\Myw��%�k�����'��8/��ja�%sȳ����N����=Y��@��.1`��H�H�$K,_K��-Z�4˶|�V����#i*+	��_���
�5�d���,�Õ����rt�j8��&�}5o����Y>��� �P��[C�g1Ҝ����Jb���4g���F�E���h��̯y��Z��*1���N���jO��=z�6��%��/
8�;Tע&���?�i��E��ևn�;��-<�TP!A�/\�55'�l��=���#�e����[D���r�_6t��ۏS�w��¹���f��O��u_�{.�Y���N3�$�=�`�T~#GL�]��	� n����>}����N�N^�[A�P��O-+]�홛[g�53��,.�ք��*���]��0�b���r�u�����zjJ�~3�p	f�=�dKY����I����i_r`y�E��P;&,- @ֈ0��������z��Zq�dks��I].]�L���yuM��L~�/2���'@Y�|�ɞ��)�I?���)��&4^Z�H�&�~�!� ���g��)�17F�*/D
0�Z���E�s�Zxa���T�d�v�M֖�#[LK&�u�8
I`O^I�3�}^��[ԗg�T\I�V�ڽ�WfSC��H���Q�ر�~���������N �>~�R0�%��k/��PQ�� h!wW�\����'x�����+�LF-�c�캋�y�]�R�^>� n�BR�I�)���Mw��~��l�B��D.�\����Uҗ��L��E���v��~�%�;vh:���h�r��w�.��`Eo.��F����=�4����Ͻ��nkc����*
)#,����8�1��wS��o�gI�00�����Ɛ�Ac�r��0�N/3�vULMK�<��Ɯ{��2�T����р�����՗��_�i\��q��ܰ�۪�:�U�ݻ#_���ay��*wF�����%���f���@ot����^� �8K�a�L���ca����:�I�����r��������b���;5�	4��Ш�Y(���O�
�F
���Y8�͝�)3�N�7﯏&���U?�����Č�@8��?	����핥��oK�Eu�ٖ���.���ѩ	t�{�6�i��:��w�"�M���	Y� ��%wrА�
d�8Ӣ��630g�5k�jY�P�U���N�J��[�Bh ��*�8�����N|��)k��`Ld-Ӧ&�G��51"Yע�g�y�Ovߙ:�7�|Y«-Lu�s��CCM{z�\�f����W6n�;.KPP�htI>L���9��)4�� y��;� �]�'PF����`h���7N�V��/�'i��ǰY����t8���°U�A:`z����|~:���M;ܩg\�*?:=
,�r�L���:3���hQS� Cwkk��ɴR�u1C �gPW��ȿ
l")7����7R3��XV�11�=��X򠍹���Wn ��o�:
���)9�'�� W�h�gY=������j�jlS6Q�q�i�<{�:�����.ֺ�#3��Da�#r!��ώ����� �P�g��躛P�e���d���[���H�{A��*��_f�Z&������)4���*��o���3�M�`�z^yGj�v��`�*�4V�M?D������Rvݕ��~Y��T}Y�J��8���&��W2;��q�؂��[GG�)����  b��}��R���g�>?L|W\'�p|��#IoG�-�ꭝ�@�O,�ǎ{���.:x�M�ߌ���Kcw��@vk�5�~<��cb��(�O��3��;�����9�ܬ�Qsg9��qG�K�i{��,N�^�TvRs�di�
�����Y� ��Di�o]u���}��z�7���i[��91w� ��)�*��P�L�@ab`6�5�0��/�)�p�>몢�MW��i��R���Z��EI�����:������8G�W�Ύ�������Dsl;[��*����߾NMI�1��< #�ɢ��B�K�ƪ��u���Ł�3e��#���i�u�Rf�s���J��\��A}��1\�?��))���ԟJ�1n%��F����Y<�>>����c��<K#�|9k��c���^�o9��Xr�ov���T|nF��&�y�b�ʤͰ���]'�{U;�� ��������i��.6~��jh�/O1<i��FF�T��8n
���LL�O�0�1*�V����n�k�q�I9���j�S����t���q�����~@@	�Ki�SUM�A�6��j�.�!���tx��xl`����_YI�Vn���l�?���&N �NT_���~ft�f����nul ��Jnu92n�l[��O�%��;߱5G.OOI��e|E��������4E���m�Ʊ\>�4�!H��N���@7L�@�QNʍ�������h�P%����Jջ�Ѧ�� ;�j��	�LA5@�c��Q�� �ZnC���U@�W�nA��AP�ȿF��j���y���RM�)Sb���y�����:-,�.m�K�󻯭>~���lh��d�]���-�w�	�tr߼ΐ��=SS3�%�ײ���j�� 0��-f����� �dې42��|*�4;����hI�QRB�d $l�%�Z��*�m�bc�fX�1��a���(:���z��W��D�� � K+�v�뿾Թr�Ԭt>����W��E�ؚ�}Ǜ��*js�C�MIN'ߞ ��v�8������ �-��b(�7E������`Jg~��c�pS����l%��.v��ɜ��� �3~&�\*g!������K�V��c.�躪]���*�8�6]�g���G��$�X��C����}���~��f�[�O6i�0m�2��΍�*��}~�ow(���J�r�#r��byj��U���p�нso�U����3�%�W����1%�z#ׄx��V���za']�_/��R����m@
��4��ހ�qV�qgO�y�;���d�!��|�� ݮi}i��P4�v��	������Q-�Ms��!h�?���lo�aUמ�tR�obb���GhoG�?ʁ\E�}��P&R���%~N�<�%��,�΄���k8���vP�ʲ��<�F���7w�Sϑ�ޔ�]�c$���M�q/��%?�L��,ʴ{#�t4�q}��.r�:�TZx8QO5���?`��!��E������#�&n]ޱ��3x%jz�p8*|�v� ���r��1��Y_O�������A\�؉H�9�dJ�i Ph<�?�n���5�R�߉R�e��0��r�ؑ��3v��k��z*螃���a�{ZľC�ߗ�f�ѐ�,M�B�v�7=�2���<?�16�1������xX�H�9��
��"�t�]]w}4s�jX�(���m��S���ܗ���E�?.��nA8�r �/�iL��׺M��]v�K�6rl�"�͟�W�����ݳ�`S��ʞ{��?\�B�����6y�4h�C�B`�� ��$<+)2kڇ�t����64��*7�Uz����U5����f��P¨�8�~ �y֊��DZL������;:$��϶ם9���r?`���U;ƀ ����Hz��X���x��R!�GR�˿������2�V�^�_�s���h��?������|�n��ZIa�<ڹq�Ӓ��βe�,=EO0���Oҥô#��[��!?F�@A���ڊ�����<�������W���Y�亜���<����p��eg����~��,��s! ^��7�����d1+�%�e�b5��Q#K�̍�w��9�C'�J�++�x�0�<�C��k�Ĉ��mE�	;����'$WL$�������Y�M����n_0ǐ�d�`Y����Ǧ|���D����>Z�QAIu�bt�>4���ٓ43�j |�J�Է� ~g!K��+Pȳ8�	�ٷPyG�%f��O��ś
���>��j:2�@���de�JuUK�ߟ�+�� L��5j`W��i��5ϒ������: c��鿤|��l�������ա�\��V��s5�0�
첆����Tĥmn�$=C7a3N�(g[�Ok(�%���O��%3�y����^���=�R�X�(�ߔ���P_�P�w��)�9�{o�|BОz�po0���uf�"�NF�W�c���/Dǎ�7�����Qp�f(f4B����M'
�ptM�n��#�i�"�����5��db�,Cr1|on��,��0�CӶ`��kD���������r#%V�ـ4H�i��XSj�2��Z�Q���Qgk����JXnN �=��R����7TĂWM�xޒ|�Z����׉�$����'s�Es�����/�j�Zb�G&?R��]���ņ��!$�[����WS],����b�t!�o3��u7���/{�--� ���}�ۻ�K��D���L�< 5�NK ��`�i}rR��e��f"��*"LC�k� ��%}���Ԍ�)|js�����G}C�����w��D9Mh�˲S�O��/��ǳ�{Е��I��,!�x91(���9'_b%�Y'x������I����/� �1P����\�G�������R�;���w�ǧa��x��o�~����999|�E5p�w�&n�I3�7W7��3߉ԅ0P`'�=�� ���pki�E@ƽu�Fj�i]IK�y���z̼cq�9����/�n�jo�ۻNF��)t}�5�=7;.p������t���*jj�����Ik�|=�DtQ�5k6x��eYU�{ۨ���x�wg(��p@�G��Zx�\�4�=q����۹e;*�.4%|ƻ�x f�� ������͓�}=���x������fj�W��!]�o�_<�H�&�y%w��D{�Oŉ��'X9u��(��a��u�
	�շ�)�"�9 g��{�Ƿ巀��>W+0�U[m+|���β�N���+ݮ�>(�퍹���������w �]Z?50��s���_^�п間�6%2��X3��R�NK�h�$9g&����VZ8��8��f^v)��pBia��)q��
��q�A+ߍw���<k�o�`�����p��r�:rE
�3{ϛh/ԗ�B}-Ӽ'�w�k�ֈ#�y�a��?ʢ'M�Ae9UG%��s��k8�B^����;�j�}ژh��v��F�!�����e��k�`�-�%M�?T��<89I���)2�Z|���J/gpX�Zu���HH'���o��J�U��83ÿ��8y�b�6���֌~v�$�V�d?-z��Ġǀ�`5:n����pҌ�!���JQ����}������M�֤6�2�m��>��@T,���PdeW3���]�,4�Js����]�'�2$�ۢ �_1Eo{3��lż�S?al�e�Tc<���D�ҍE��!BI���,�=�����)�V�2�go�QEyo���VX����f���x���	����?����@��M�:���ۤ"�O�-��R�r�e_"���sD�f4�#�q�m��1����w\5���|�i�V�gR#@��=~�{z#W���w���A�"P8��"#�_fD+��α��I��&�	�uM#��ݏ�v �:0���٬qeWMsiGX'2�<k�}�J���Xx��~l�}#�Tʢ3K�$M�OR�G&��:@���3�^6 ��gՋᤳ+���R�C��-�2���(������-]�O�_���X��Շ�*��(��NW�= �p��������GcIzn�`ߥ|�d�ூ�R/H�S���N#���?ؗ�o�2G���&Kw
�d��Y�L�+ʄ��_�w�V���J�w���[�_*�C� �w�]A�b�*����P�9�+I �1_�j��5�A_%�(|,3��c�����mB�n�پVx��G8�%�l0�%��.FT��KQ�<�/�:��^���{EJ*��eʻr���g"!��p`����D�o���h�A�e�\��t������qh^z?b��������m������5rZ�u����m��C���b��/������v�������[r��P�����ucD��`hO�S	.��}O���R�"�?�ӊ�m�"F��?1=I����~�J̪	r���}����˾����Ajb��β���O��a9Z�lq��źCZ�za9&�[�.�]��ݍ_��! Q�fs��z}Ҽ�+|Hz��
�L�����"�k&�j�q������z�F!+"N�fQ~v-���2���F��k
�0�����2��(�tWg.;4o_�)`I� ��t�8�� '�o϶�L~�;1_0�<p��.�!^�W�Ԧ�'����
��K���MH��]3z��ă��?/�vؿ��UM�ƻ�<���q�t�}�Ef#����u7ߨ�Z����dZ�e�V�H�[���7�k��|"��T3�k6]ɉ\�K#��Wd�g�{�5S:�͊ ��K�&�~�rb1Kc
]2_0H �%��}���\��p)���m9n�{��0.cqcGk��RP ��M�҃{�iP7�"�Wcؼ�Do�sL�@<}j�q̉�O��H_�n�)��e��E���Y�Ŏ� �Ќ�	�衏���I�7n|�%n.�К
��Ȑm	�Y4x�R6�����T�,�F�f��Q�[!lz`H���]$f����J��p�D�W��������ty����7m��ԧ_��"v�挌�;7�N�L1��. p+JT���q'm7\b�񟳜
/��z�j���_2���O��������0[4�z������KYG����������&���ip�O�p s�Ǒ�|*���n+"x�f��{�Ǣ�no)��je�x�T��.T5�a�~�����$(�[#�
�ۅ�>�xܒ�MJJĹ�C���A��!����A4?e�G�-n�*ׂ�r<8
 W߃���0y� 8�O��ח�8܏"�j ��U�Ź��py���N�JE)��[��<|�O��K���
LL 
���I��w�Em��W�3� �Xqck��I��
(A���ik�[���w�x���2�RW2�ޣ��ez�8���6n%�Č>B�qJOb8O��8i��yT�";F	qn����o&�M��#JI݅:�Y�1�J�e���x ?:n�ʎ���,���ƞ��h�f�O�oߊI,�/n{c��v-D��Õ����KK+g�#�߸�r�p�#�b�he#����ǅ������a��Dv	I���!FR~$��K�.��m����u����:���S=\]�p^e�oА�|�wX͈[4]�a'��Ɉ�8�-�T��a��<�j�g��XY���#�k�q�.�����Y֜�׎�O���;C�d����^7���H~E(t��Iv��M�6�Y�9��$+����ƀO�Y���n4S�@�����J��w��:�|�V���$3s��`��$7#��g�E�?0�G�9�W���̱]T�o�mx�8W_̉kI	�V|�  �����	�>���{��n�{�J�D��ZQi���O3�u�Uu&G �7P��Vּ��ޭ���n���-F�n��k��c����%���5�	|��XB��!���7�u8.��ő�@E_>O�S.x�FB!5 ������S��ZQ�Q1��|�S����;��s�O�p�x���lƨw6�#\�*~�;,06^�9��ɱ�:���@�8����!�s��Ј�$W �#���try"�A6�5��{<����E�\�?�GiFZ�	���2uuM�)P�ҿ����l���0հ��Va%�{���c�lߗ���I-}�U����� �w�k����NA ?��>M�Ep� ����D׫���u�j��xtl��m=짒�������p�Yx�ߌt���,F��� GR.�[�������}�gL���"�o�E`_����m�����n��$ƍ' �잒�ړ�R�m�(�@�
4Q�N��ſO�כb�ɒƁ�?W(@9o5̈�� �`<�i���o_�G"��G��08���"��C�.-c6����J�� �%�V@��?3(a���a��Gs� ������)@�?/�w��K����6����]r��v���܉���ޞu�b���$7��;@�t������������Pݜ9p���Θ&�` #�]��SS�LB-��એ���Y�l���V�O:N�������#fS�c_*72u¬���Ǯ��<z�4N�H���g88�*��=�2�O�����5U�ߋp�;�/G����o^#CK�Zas;�I�nG���=+���7#�d�ĉK�@��������<��6�̅i�TD=^
�J�7ˌ�����4�m��5Q�4�r�W��"͆ђ��8@{t���	��R9}� ������?�O�ɀ&�"�]8���\\�6��ϐy�;@b���om�7�p�w�ڪ��Ȳ��'!�#s�����9t`�,v��K:^T��4���d��J� �u�������S�#W
�/
؅�-�\���$c�^��]����Z���'٨��^���w^9n���M[[?�/�E����%��Fo����`1w�.��,�H�(����� `��x�ŝw�D���G�lJ�h�7�"��XW���^Q%��^?�7���a'D`_)��sA���̂�\\ o��m�}RВ��B}�x(��`�426���*X�K���F3h�_�B{Ė� ~,O��N&^���j�z�ǆa�g�֫�9�~��oٺ�v*>1�p�14�����{d��t��ut�8s+?k��p�� �*���(��0E�L����f�i��LĝM��ȹ�����o�d H��B(�����)�ܒ���Lj� Jp�uO&'SJ[����Uu�^�O���>��qL�Sm�	�Գ_؉Ђ��!-�vü7v�< �K�W�d�U��NZ2<B+ce
F�a���B��t�ZZzI�qG�8��=%���1N8�9�EUDj�t>P[T��������K:z�i$�dh,J�>��yS����<K�� ���)�%�C�>ޤha�7F��*�үx�s"�yf{�Jյ��G
�����|�I�����g/(�5��i؋���.��$|�W�?Ĥ�x432�� �X�s�X���V@J� ���e��a;���zv9��$��bu�ˎ��1n�Vd�I��D�s;�Nю`�$�LXE�I]1*/]��6�R<���Y}��-y������g���d�^�4�����ǳ���H��BW���pj�D��y�{n<K�Qꀈq�Q�����#����@3�b6�H���p����p�X��!I�K���NW�2[�����-�I���"�?L�Bt���޼��h��IӞZ�Z��cR@g��C�[�� A���h�7�-�uv=�����$]ЙGih��ߚUN�����63'7���~ْ��[�uVo ��"Ыn�B��Ϲ������I��	^��RS����4�?�P,ႏ��rk�!rk��E�uW�݉�l�%�!���ͦ�����"��5��6���`� �s����j�}f��[��C�W��5
�����,��HY�M)����,�|c�h�%�����ϖ�!�?#L�Y��BU��$�6=�Cw�.���v�'�O'�t���p"+E�E���LRi���4�ӽ���Ռ��(1e�]��M�`�0�3�FXuTTOǾ�^��g4S�|��KWB��]���U����8��p�|�ڗ7��$�D;ht{����=r����:\��AG�]�9D��v^!pE��t��*�r/P+�HV�����G\!+nX���?"J�.�ˏ����KOL�e�κ%��
��qy�&q��A�J������o�ʾ5Y}v�W����J�<�\�cｚ��8;2�Y��L�B,b�q@�Q
�ӱ�[p~�Wxˊ,�!)�:����U89O�8X��VK�ߤ��?|����W
)�#
[�6��F�$�V�M?�\=�kh4A����Г/� ������S��^�q*�	���@��3���:[���Θv�D��o%��$��� ������>�E�ȇt�N����2�8R"y�-κ�B$B����n�z�n�YOv$z5M(+�靥r�{�ě���Plxv�&t��uaGx�鄂�V���0�_0�Bi P�'r��`j@��s�3���/:����uN,K;���	Y}��R8���U!�$��"SUo%J�~���aоvw�@��Q�D0H�^�׊�'�(��V�a���0<�LH�k�Aχ�x6��:>p���[��tM��e�S�	�u����W�Bm�c�5FII2B�UAaL�}	��n��<���o�W% <��K�1#�<!�w-�{ �^M��$�x�e���4Hj�m��L�^xZJ�^�)C�(q�Ռ���*7A�$��"-����4@\�W<�V�m1�)�?UE@�ݘam�{1�J��Hvm-�|�_�0 �qc�S��o"�ħ����HJU[Q���=`h��д�G�mg�h�u ���ܚ�U�gg��í���(��ek������n$�D��i7�3���E8`ht�J�M�9M��v��+��|%n��$o���|I��$9p'}$� $wX�V7����~T/�~��F�CY���*�c���:W��!��t:ŭ�_C���S� j!�C�a��3㮶O�$b@L��a��4�|�$DM�n�->;\��6d|q����^�/bhp��U����?��t�����u{;�3K�⼼��K�.k3+�qA�M"��z>�Ufi����ű�J!�R��ᅌ��/�Mk��"�F��E�-�����U����+�#�w�F�Δ{�[�]�洒p�`�[��O�{+]i`�q�J_�.�L{���:�{�=	��O���R��wl���乶�x$�:���:��������2�������~T_��9#*	�a�}�ʽ9ߗ��4��u�¦>'�)�kx�7?�5n�e��W1��g��֪��y��;Ny���"_�vHq�����޹b�H� ��'Ǭ�ܲST��TZ�;�9�<���q�*��4d?��������a�M��L��M}�~��o��Ԩ�l��M9;�ס����U�g�;m����b�Y�^5����;bs���,�#g�فF>���&'��b%�rn''���\�;�Å�]�|�R�媼�]��u�ɓtĤ�[L��u������~�^��M���C�h%�ҳ0s^�E=��gDy�<P�ܭ����D��ٹ�F�6���F�:F���gE�K�x%Cϛ�� %'�5�n�_���1V
�������q�L�Wʀ���z���UJ�w1?��C��<�o'K��w�D�v��(#:Z^��I&F=��6}�V}���'-=��R:xK�K(���2�����@�U�	����f{ ��R͙jD�IG`�m�OG�4�0��.Y���������~!��.5@��8j�Y1]�>8��C�t-����ɍ>� 0��̀cG��d�Q�dr�f�']6�
�|��c@A���!�_�y�����q�HY�Ye�[�ͮO�;[?�L����%!�����w�t�nY�g]B�A�y�'M�a�j�^g��5\J��Ԇ��l��=N��X`ή����	m����
�3k]�
_V���!-��P̈c�濜�F���Z������Ţ�-���䆎���_��/%͢����oA�Ք �ٳħ� �X�F߮�HgkB[*R� �َ��j�`^k��!��^맹����T"��p��j��uJ�&���;��oS�d	߁��x�M)��[�!��N���e�7[��;��x�<���XZ����V/��BdѴb`�#�F\В��E�8��y����a��W�T�a�mZ��Z�
e=���u�m���t�����ɏ�|������Շ����vMծ�����a��p 5�Z�M�����܊2"�B���a�	E�0����p����qf��ɀ�w�0�*��c�mu�[���j��7nK>zv6&'���N��!���˒�Uxk����QB�bz�����2#�{���x���o�hMp�A�����b��,�@��D���(��1��\Ǣ�S��� i�C�L�^�5��'�4�q���V�Gx=��5����ݎÞl�܄���3N����8���m���eb<�����&sr$��.}��}G��T�)>�I��N��|]\\���k-��+��9�1�W�=�	{ڹ�
�ˮyoQ:5�B�Բp��K�!���v�9��k�p��લ�G�#跔ä���M����Z;�4�Z����ܪ���"���?�����L� ��)/��|�����I���Sy��ʧ�m���N����A!��ׁ��|a_)��>�t�ǲ�}'3Β@#z?N����l�)W�׍��D�8A�ژ�3����D�\`����²]�Ct�����绡��@�\���9n�&�X���UUU%n���Aw�u�PtgB�@YZ>MȈ��t<��N�J���ɨ{�]���0S
�p��͏�����/�F�6������(oi.�}� ��-=����|L�g	���8�_��n"�v�e��V[i��z�v&�;�g��T�?�ZF��b�^2�i�T��뾻!b~(��P.'��v�8�b���̴h��c�Ryا���G�ג���9���(��y�	s��C��.u&�[}�+��=�Ib8��C���*�`�w=xg�a�QMp�Ó�%u��n�$Vr�����3����IPI�p��i�{�z�5|=�h%0a��{eb�]�o q���܄-����ҽ��ݨ�h�Z 76�$i�N̿�è9�xG;�X#���!��q�.�zǴ�R1/�i��<�2��ry�������}=⾂-G������lKD�1�9�!������d�?�2A[�"�������%j���ڄ%�^o�_�l*�_o�+l]QA���:�˿Jpo��%����������o�C�އ^����%�ϋw��YJn�#
#p�9��:
��.,�J�Q;�&$�a8Wn�]��$��$WI�:7�����o6� ���J�7��W<�z���ބ�`���/�E�2���_#F�������Ozfu+}�-��"�M��,vk�����0m[���sa=�� Jw��`����J�u���t���Bo�ǮU۞+�	�F�O���0]Xp����~EI���l���_\{PN�i>w�������uZV�%�=���j�y�Vn���t���#Z�C�6(x��C�YO�&�R]��*��s�F=��mG��۱U^u�\w-�m����� G��g���X����K�(���d%4����3ٷ�s�@�%�+�)�mCj � ��4��F�t&�H�#;����5��Ꝯ�enl�k���d�1C�d��+M�A�n��V�u�p$���Q~�f��F<$]�}��2�*��b�#�>�����7����#C��~,�L�d�D]<7u9����˿M�7.��9��þ	��B�}v����O;���g)^��Dj�Ğ>����營��մ<�4�V�UEnG��`_/�G�����_&0g�85�P��Y��K��@�e�~+���=�sږ!բ�t'}�q}T�|.7��!'-O�lLA:��O��.����8�x��n�bW<Y�~ٳ���иQLZ����H��i�K箩�ܭs�҂t;&X�f}�;AR�ŞN����B��
�B�:�X�i�Ń~P��c�+� U=n-x��b�xF��<ΡR`�{���I��Nʂ�A7���l��/N��P6�m�c�������D{���1�L�L��p/㼓�+�����-U_-^n^a�gE���T��C����L�n�č�>dm�-�K(�$�|�70?N�9��&��]�dϽ��,'��M�b�#�n�3���m%�7l��'
o�b
���=��m�ⱑ��ɹ?f���)��@R-�~D�g��S���J��g��"�1���8O ��{'A��wn�Ћ�Ԑj(��DJ�z�Ԟj4/�&��g������]#w>������ ��C�9~0f�1�sI;����M�ޡ���9��K2|��[�A�]���6���;�ş�q��w��#S�N�zB�Ͷ�!Eɼ��+�	��#=x�̟�o����K��h����Im _�K}�.����4��11��{J�>�].֎�u�w9�z�x�x�؞z�`��S�e�ޟ_��N������[kb������}'P���v�ؒi{����F��g�o�Ǥi�j��-W�Ӗ��}%܍���$�\}�]?������W�PT�L������I�/%�dhudv^�D�Lې=z�Åŕ��~V��Ы����W��:8���:�����GE���M{�x�^�d5y���ǳ����Ά�z���X�Cp2���C��ҕ�bG4o?��C벬=��Kt��[5����u��ۻx�e��������z|�>�״�>��H|k�߳V���v��Ѯ
)������o��q�����;L�&���6��\(h��y5391�p���w1wڻ��6��zj�T�@�&bCӽ��,@p��\���$%����� R�/z|}W�)����m�nh!F���6ɴ6-�ӓ瑩��ܶ��RMM(����4����fsuhOY����=L
V��� Z[�U`��Da���q�P��|�k}�.jw�݉Ι)�8����RQ�st)쓗m^���8�1N������L�M݈f����[�6�ɭsڄ=�� x��7�����W<�s���}���!�:�
?\�?W��2�~%Q��O�G��~S�fڂA1O�b����+���XUf�l���ٯ����X��3�q3��pY~�
|�x}G��6)�QF�ӂIb�ʀ�{	�9
�"��=�H�{c<
F��� �E1����?���z(8��\�v��|)���d�KgR���@�#)o�9Q�VT49	x�(�����έ���ic���Bu ,� ��ߘ���Q���`����"��n���N|�U��c�w�z�TpHtVW��R[\v�f�?���u���%2
�|��, m�ω�.��u�F���Κ�{0��u#��+���:���l,/׭t{��[/�KᅇLN���L=)���i����`��S��A����c�o*z�ĭ��� �r�6r��Y0���'����dk����3�����S_���;�t�t) �ݩtwJww�(� �Jw7���]Cw�;�}���e�Y�}���9��Ĝ�������e��:wJ��b�W��Iv�ӣ������a�8��f����y#&� �^Z}��b�M��|��SҼJ����ڣ���%���&fDV�CDֱ^����rsE�ͪBa�MHi�܇6�(m��^��v+�fQ����u�󔃩uB��	_�h��y,]����8��D�-ЖuVh���4����U9�5+�m�&?b=�.$G�BqF]\ę�{���]{\���z!�C�����"��� dw����r5��b2Yy�b��oK|NN��TAc����[X��#R�5���⏞���(8� 2j��	|.j�I�&����C��~��q���6�S�]N�ǭ�0�Ex����b�A(&�Æ���M�����G���u�����p-]�1�[u~䀣Ⱥ��p������M�z�a��G2Q����);!���qr�I����"��n�:�V��c�֭�[�s�Z^�N�V'U"������IQ��� T��-G�#w����Xa����0(�g�^��l�+rw��$BB�l}3`���(��\xg�pR\�Qͅ�<�@�'�?$�/���q�M6��`�KHRۭB��:���d3}Hk񥀄g�P����8�������3p+��������7��]s㒚��h@�ɓ�~�&��=1~[Xg?צf���@/E@���0��F9\,���Zϫ��8T��'����i�/c/".<>v�ݧ
P�=׳Pv��&��;���v�[�i�X�`؟��L�K:�~@��_�b��.�ML����^��T��,��V0U��v� �%��\�5��Ȕ��3�����pk���E�t�c�ܬ)UZƏ|T��ˁ��%�����P`XY�{���K;�e��:/7ӆ/�H�Y�;~N�o+��,eU��6!'OrՂ�����]V�A��V�U��G7ux��O�������I�w;;w"m�ߠ�]zF�͉���u(��U�U@a*�10�l�� Ph|����ͅ����t-=���ЏU+�xE�D"�K�,v�%pK�>߬��o�̡��_#B�2�\C�i8���0�%z�sB+�ؤ�OV����D�2�\E�5���3�a�Uϰ�$��t�9�H@3�� !�4�[ѯ�߈/�N��S�D�Ҋ��\�(����_EO|�C������mk�b�,�ԁ���M"$��`\`�gO�b��|ء<�dL�����y��$:Fo����z��|k|� �>��Y.�1
�#T�ʖ~me�3��p��HcH�bG�_X�ّ��"4��=��C`f >��V����泹*�eNd8��Ƨ5>-ZV�]C6�N+��TI�;�lMU�|�~2�qy5�Qd���N���J�!�ey�"�' -�	��dM*	��Pؘv�0����
��)Dw-�O1��5 �#RA�ǝ�u����g/uw�J�p�h�G��Vw�/�[����:�<�$�~�����4_3� ����v�@����C�����%ص���[����v�z{�}�)\��y�p��{��U��?���� ���Zh��Ρ ��l�J�\�D<�Sa)Ja���2(��L΋���Q��������t����?ɑ�W�ܢ��fz�"u�����r�"����ԕ�h&�L
Raq�g��2�cSj����r�+<p�<h`����4]̳�[d�򄞎��:��� ����-;|�E�,�]��%�ÖPۈ7	s{
���h��q�smp�ݰ�Y@
���?Y-\}�r1��XW�碅�v�9�s��!�7K-vF����[A�d� ��o�{W��q��C�?�Xq��k^�w����pRߏ���+�����K�g�q±2�-Z><h>����ڨ�4�`��b��B5>^Y���p��w��oS��ntə6	���^�p�{ި���8ɴ/'����f����M��/f�L�b���qX_��;���>F���%2�y���$�$s?�c�}@�7�7*�6��+;ݖo���+f�|
�N�4�mč�@k	���G�<R=����Ӎpۇv��@��.���Kj���1��w��N���:��o5�>Y��s__�j9�=�55^N4v5�5�{���35K���h%:s���Sr/ 3?�j��SO�<}V.f�B��U>��/�N&Gn�]�묦�f�e.���o���x�`W�$V~G��3.�䎮�^-��k�Pa���Y�߅��k�	�	��G��h�~��̎Ku�-~N@�p����ՏVW�Z3��'���",�;>t�A΃��I�ך�ko�����iM���qPf�߸��E�sc9"F\@vO[�A�o��H}�dH�[�^8���倛�ϭy �����,�*����]}��a����W��64x�4B�(�>��6���w�J�A=������������jW^���3�Mt��o�� q�(KH������h�P��4<��`��t�֣ ��~O�O����0��P�sF��AL���y�&���"��-��'���f(�S���D�"��g)�W��
q̓+��\V5�=��w�M�R�T��Ӿ|��>�WW&�+Df��������|�64�� ��D@`y�����Ύ�_^��AW������`��g��TG�����e��/`���E�I$�a6"rk�r���J�pj	v[!��8��&|F:�n�ԄO3V0�I,�+��mUV���W�������^���9 !���:4xN����WR����c�z���V�{�q���}$��7Oʑ�)�$��+�n�l�3�w�d=I�0#���-�Ѩ�F
8PJ��?z �9gb�[�z���)E�+�����x�'�����7���@yl�S�E#�~����dIk_F��=9�K�f���
�#Xd�$����e���S����:s�d�@��X\�g�y�Ƕ��2&�^�f�\��x�7w���X�W�,�8�B	�\��HIIMܯ^�x'�@wW\|j\b�y�ZO!�sͤ����$U��Z�+D�'���־j��k���D�FQ6����Q�0\I˾ծd"Y�fsv����ڗ`��KZ ��z��΋X��QHW�Y@�dն�a ��Ĝ) �V��
�F�˳��ᨐo�jԗ�+$ɦd��S��`���=�"y�.i7A��5\ae��:�/'�x�ǁ��NT)8I.2�������~n���b�UfPwG�+S��V�I�=����q5�셻���HW�7樎6ׯ�;�#�˔g+�ˮ��J%�d{�h�d�fQ�����%�&$�ߟ{T��������O���=�"���ub+!������rf�GZbn5�8_��>�`��i��D|���`�zo��-�[P���cZ)��;ɨ~����#*��y�kL�.�����8�!Q��J?�l�H����B����?�)�N���gW�ѣh!�vQbs��8������Y�LB�1,"�p��V��Z�A�9I����4�	��9|ʬ�z6=r�Y����_����I6���r��[��r�6��
Z��kR(;��c��Sc���ᲃ6%H����S�F�y���ڂI���X���݁�-:�P�&z	^�%�Ђ<�S����C|�u���OЧ�3���M�����ء�)'O�'��-q�k���r�MR�����w��̛:mw� ��^�m�Y���x�����?�n��h���\�ߨӠK�J�����w�U��
-C���CF�a�FX�$�����jA�}Y���D�6�ۤ��Y.ӼS��S�K�/�{�R��ѫ6��s���C���"x����H�B��m,5�F�^�������w:�A��{ǳLX r�aA�ݩ5l��/��]e ��?\�hBb�ˁ����?*�W��Կ:SQ�.�O�W_�d��! p�˹
�i�8�ەZ����N�B��%k9��Yr�Ɏ+_#����BG+�/�+�����������ٷ�S���lĹ�!�5}R2����-���!���>,	�h�W�	w�W�Sx�<苬�6��V�?����Gm�v7[A����^��>@^*���|!q�$Z�O]ݢ�u55����Ī�L�T��ԟ�큟?���-�h�pj�"��7=z�9�nO1��,�`�s'�t�����������J^�� 0)&nh��^�'8�S,'�%̭~=��.9�J=�G����}P����{�F�?������B�ٻh<��|�^^n��;�������I#\N>�.d|67<���+�o��ب�������v7�*�����ub���5_�Io�޻Ce�u�i% ^@B�hto1�C���_mQ���ߜʾ� `#��ДCޙBt�ݭu�>�&Z。`y�,̕`g�7X$��y����"O�/��/��46��$��I�t���n�FfVwĺ"�7�C3��A��M�T��2M�ӳWЮ�m܁4-�6��I�u$��^��)�eNnn��#{�������꽕����h47wwkOO-P�Rj@��6j}���l@����4�B^�\��$��`���D�;���HY6�-g�W�����<�x�9sɍ�\4���������yf	)^�>�?y�&�̾\fG���wL]�ႎ�2>�_��z8�
�Z�@(��rEee��V�ia����>�U�r �l��]C's'�>U��mI��o�k?S-�w{<�p�|�W���K�ٮ�Ѐ}d[�^i���M"W�6� }�%W+!�m�|0�����U!xf>`9�q
P��&N��~yRZ��㔏팠D��y���/7$��1�^��2~U?`���������#��{2R�l�'Qb�g�5�%���������f́t��d__x41o�x/��2yӎ�{��"`�1�,Z�ӄn�0�8�͐�	+|����y�k�|y�;���g��qI����}b��UxƲg������]giw�ԧ�F���a:l��ڦ�ǉ��p8E���W95�hSsa����%�����_�-6}6Xv��~y�Ys�������+������������zjeb"��e�rg(	:����v�8e�����aU�x�I3BB�;�	�_��L?>ko�q��'0���o��b�I�>Y��E��vF
q�{�ǻ7�S�R[E!;��D@���!r3��ى�<�]5������v�R�u����y��0���ʝ/�w�sZI��c�s]��G�9~�6������D�PF2ϛ����G��Q�"A~řv	j�#�"?��Q�<P����%{��������L����^{̀)4Hn)B�P��b9��wCO�ThjBDȯ� (V������ynڸ�m��1��,,g)���8�ԷP�6�:��m��T�����j,N:*��(���q^<�X���s��f$�޷$^�	7���6�����`j�x��e����
)G,+vr��q]lzf�@(S��|��*��������EzP����ې��?�	��R~�c��P�F�nb�2��K&,?\�tQ����=�j��4��"-�w9��g�i~p�*����q/7w4W9/-����@C���΋/R�U����m���m��,<���J�T���|ʊ#��$�흔q� �\m|���с����sF��9+n(;Si��Sْ_�Pa���Ɩ�c��QAz��3C�+-�/c��Ȋ��_-O�x�Ϧ��+h��q��:	y�㈀S���Z7���/� ������]M��e����W4�>��d^����U�O�+1@�E�{�ΏI;"R�/e2�Ww/��@�Av�vu@Ӂ�ׅ���?�l�מ��Yj6��aR�ɳn�<�+�/~w��S4OCC��~7�Gz%W�Lzz��
�}{�()6��/���%����7r6m�;��+��CjɳH�ܜ�NQt9s��+O?� ���^����y|��E��T�̇��� w/ZiiH
/ʣ��eM|��z�t
�kc��O����e|��[�����" &�H�Ñ�;�I���$�6:z��;�t�m�����3O`4�B�-w�o����G6'�����胡{��^���v����Z(����ȶ:``�:�����cp���zC����x�e����8\v�����G�`����-�|�E٣�E>%��ĽG�S�^:F����nƔb���;h��L4Z�c���iɃ�r��P����'F��>D�01��R#��G��M��Y".[�=4P��:'�t����J����hQ�g"�=��:�M��Op7{d��yJ�قG�f3���J��k��a���^H�=��	I�*؞���tv~j�ȶ��_#��/��k�v�|lE���meaHZ)�&S�����1�(���c�|�;�x��^���,�r��]����W ,��4��khSa�͎f������aڋ�����������bR�n�6Q Lצl�n�%���{�H0Yz�^`pI\ ߴ� \�B��<�v@���RP2��*]g3?a� ә�i��w�K?=n���@�)LZQb��dl�9.Q�J�m�[�в?�UXJ�Z�Z������o�v�������M'��μc�S�(��@h��Ɖ	F�J�������i�|�x�5�������@
��1
̼-�u�&�
7j��p�e*t� $��q��ݤ�v�ޯ��)�Jm� {J�c����:]aRŃ�0ݫ��*�l�%_����Stm|�f�g#�O0A��`�Ō��_-�r�w.�u1�T��[�a\���O*~�::*� T<��`�K���Z�֮C���YrI׸q;���$��ġ�|�,�e�I�����f�[�U�C�<�����i�6��{����Yޟ�_W/�!��@(�V�xzO�v��� V�?w5�-�pS��&{&�	G9��f�<8EE�1�h�g���y*�_Prfz�D�����|�j\׷88ʓ��
�M���#u�W���m��̶HYHd6,mp٭<�v���7K�:��֩�N���ԝ����hO{�j�;�KY�ߨ�>�)���+�9}L�e�rS��~j�&�V���#�L
�}0y��O�]�ǖ��H.��[����p��Y������u��j���k�q��Q���d�͋�t��uM�`:�����ǠC��7d �pOX��bF�ꕦ�P�* �q6d}�D�i��t��Lɉ�cc?�Z�JZ��&�2䨁� ܎d�U�2[�����O^�{b�M)�[�U�3ik!,0��/�*oS��_�c���9�@�Տ��2K�S�u͗,���5���=�k����:&\G6����}�.^�q7�(b$9�D��j�s2�UW�M�����~.9�OO��?�n�8��Tk���%S󒯂4��Ij����<��84UI��X������S!@A�/��c���֞�J��N�zϦ�nl�G���\�m�P���憺��� ��d�8�4Y5U}K��id�c��n�#�R�m�t?�*��a��S��wfU���� �+�S���<����ܒ��ն���;=�!�=I�/'&� s7y�#vgr����c��(�!�n����'�����͢�m��enɕ�� ���k�0?��>�h���G�ݕ�6<I%$�)ô��{������r_�Po:XٕG�*q5KV�o<���^��acWW���倛qz5��'�f�uw��«0�C�T�Wi��
��e ��g>(��<�]�~M8��tk���pW��~�z��X��ԑ�ۖW9t�2h
10[H�����Va7C��Ҍ����w�V.k.�n�њ]�>#��� �o�ht��S�㶦罖.\���V������x��'1�0$v��:aA4��V7��6�.15�����Y4ǳLx�@8��fKvO�a���=��~�Ă��P`���ƶ�;�%p�����1��b�<��~���u�j��e���@�b��&Õ���ayw����\T\<d�Ze�Q��[��-��e��,�Y�褱�Z��t|�L?w{P�5�ŝ�[8̡��fR���ت.&y,�����|��E�s��Q9��\uVח5=��xfqcyϘ$�H����i��nu�D�H6���q��`��[S�s���=C���f�Z��BX��ˆ��z\���eOd
yc�)�u?/���rZ!��!�2.<��Z������5��Z�����V��.��^�v��p�wܖSIN�K��/m�@�|�����x:�*�F��a
����k����y~3Ȅ�4����� ���P.��-6�������NWoY,�ؼ��W6@Ew�I�m_+>&��i�4�
�]�=�i��#��*���jD�,[�50`bFJ�E�SS{�����E5v�\P��I\5�g��ϩm&����gǄ��q�#{�]�u�hJ�l}����f���cc�"rl���>��������C`&qL�~:l�'zM`/7**��m��~Ӆk�����+�1;̰ fM��n�{d��C[E��i�1�I@/4�l��@��*�B�vh!�,~	ꃄK�^�t��d���������w��"���/��sf����.�����	�S�4|�n�;��{9���F5�o��ֱ�bY����.b��d�jI/ \��7���*l�Y��.���	V�"�3�+rI�48����_?�|����ii�Zf��ߊ�/���exkS� CZ��h���ڡD{Cň�j��z>���FÝ�������n�d�_Y��ҟX��1��ݫ*yԮc�v�AJպ�>nNK��#����ba��{7}�|��p_W�BG���uW1%$th�$�1�̜�����C�jT�i(�+��%fK��ww�u�)S�76~<Yi��Ì��y}
;�tZQY�p"���[Ѿ=�ss}���\�74d����7���iI�Bh9�S8��'�56�E$�=Nb�j$4�}Ӯ��Spc���b���O�keT���ǟ�`�����x��"(|�l)���9x�b�/J@�c�=���-�*����W@��%��;LL�iX�����zzz���Pu����O7��ON���V�+��P�؎^�_[��+0�?&֚����O�!X�ؘ���iE��Ki��h�tH3|\�M1]O����%�ld�U0x�ǅ���cz����w����Ǚ��D�\���W6����\gܻ�o�ps�Π��/}>V�gV�-9l
Ρ)3�	c�g7�L�xk;����vA�3e�DII���>�@����p�7.n�HӨ����7]�M���)0��`ʥ/�����$.۶O5D#&s��V�U&������ɖM�Kx88	��`�ε�f����(j���L�o�*7Tg:L\��O�~0�o;��_��t^�u$�!�9Y E5F�a��`�O2�\ �t6ѣQ�0w�+��S���kݻY*3#��p������_�,k
6��|����Z&�<||t�7�t�L Lundz�����I�� �/;1]�c���s��͏�x�Iتd㻱H�}^J�2I:���� 
�RE쭲�U�����=}w��,��D�z�� �B�D��^.�s`�(�� ��naG���%B�LZ<�/��e��yl��5�A���G��`��������!\\ p��-�(��\8y�}PP����\[�0
<Lxxu_���{�J��C����_ēK�������.�V�U�}LN�|�Q���:���.w�Hھx����6��2��B&L�I�ѧF?�h"���΀|������@S)xk@.��t�^�|6N����oK���}Ǚ|�]����b�ư(9��EM���#����B.O8��R$8#�<(�}ӚCBG�Α�QS}||�s0<Zj����>G��N���� ��3����*��d�z:�����H~����L�03�oqos 1�U�&�lE�ŵ׎\��{E$�솆0\O|�o=]�O���Ō�N.KR*;J	�?JV,�U��kB8Rb`.�c�W���(�&f����j�&
u��	
L���l�_l��E����h�`ʬ�`�oH����M��&�);��A �M �G�.΄""��'��w���ט/;<��M�Ar��R3�<p�������?-X0.EF주m���,�%�j����{{��N1�>]3R�W��������h� �$�64�x�/�	t��%�>��C~̹?�$� TJ�/dX�:��4)�_�����J�+_x����cL�YXX���Z��u�&�zb~K>���;N~������.�J�y��C`���ֺ}X=/�[�]�ޑ��������C ���X������W��<?Z��R��6J��ʐ]���.)\
���w��R I+�^��@��,��E0��D0P��k5���Jk�I�8:�(���K�7y[�x ս:ƇTS��sh(���333�4M�W>��S�&e�AnU��a3��y-5�i�Aie'8��'�T��Аtܾj��
cy::T�د�Q�>�#���E��ix[��z��)y����P��N�X}G��L�~������+:�B�ŶЉ��O���=P/=�k��W������j�`4Pv�HC0��o���"����HQ˒�cab*3���璧,�܀��R�~��-.�˃u��%��) ���.C}�C����C���\mF�K³�w��բ*������-�R��Y��T�X5����� d#�$��&�ɿ�pQ1z{��FQ��U�7t��k�CRMA�R��nZ�f��ޠ�`� `2o=����uc	|`�x<90�=1�I�0�t���{���
y�,2#�+�x�X��w�[r��G���stt4V�H�v�@E�����iT W.d����hs�5����|�=#���K�o؛`�a���\F��K+d􆃣�;��10�?�=�Q҃i��ܗ��Y�B����4�d50d��Plrd�l4_$	��{�>�Q�o,NO�!���o~����q$$*�F��\����c|��A�`����)Ea����6�=^tt��l�8X"�o����#�5�����^�}��h~פx��'�X>SS������ތ�O{I(}�K�%��A����ȆFz�P�����y�y�v�f���[Cf)_P���(�(�N��
*PC�HEʵ/~s(Ja�O��c��D�1�[o��ZH����E�E�%��zA�W %�����q:�������k�,3���#��������g��΢N>�*�8��L>�����[Z�A�j�ù��o�ͮ���]6SJ�|�Yxr�B�1�J�L�Ҥ�������;9d�߱@�@���������J��|Q�<��H�J 8��b���Y��U�7�{��No�K�_�I�������{��BH�\ۄu>�������F���F���s1�Յ���r,����a<��V���ʇ��  �����<�Z���[���4�j�&����\-9/�t�`{dx[{=�1�~��6ۨ� _ܖH�[���^L@b�G�)�z:�гh{	��|�Ҟ ~���9�~����'�7���bb�%�k@�ɿ�x_���h������3^��>gz��1����/O��[�;G-��j��z��RRʵ��,d���=�!/wdS>��J�E̲w�P�ٍF'��Ԃ�k#�_��&��ZW~6��f��g��ѕ��6B1���uo�R��0+A�GY �B����Ub�P��<���эA��T��ݎ���P�g�<K����b�r�...-��}ww7-=��ɰ%Gve�����Nyy�VIIɋOUMMhz:	11q|@��d���������$�H���+��,(�3bx�
�]ͻu�ea��M����e�M����.�>&��WCC��mnlDR���
�����~}�Xgw"����0!YHd���/,�C��i���0{�� �R����T��ґp�M x �B1��[Q��koR�;7c><Xz,�Cc��6�Ɂ,�U� 
�_�o�ۀ8=udr~���SP	p��b>����RPPptw�\TDd����|�����<[��( iT��TnR)'9�U�:�r@?�C���-m����qY]�;ZZ��[ma
��3k/n�j2�����5�;l��Q��E�G�����H�÷����a
w��D0�smK�N"�u�XN��f��5� K��@%����B<PIٷql�9�������9��k�C�k�&���5�	��� �t�м��5�sj����x�5�R_QVV�ښnbr2���!u��e��А�=wD��T�&���f��f"2���hй&�U�֔=�9*���k�s���y�B
��0�7]��(o򧧋ۭ�`��z}�^����q��'�[�Sq��x�K���Fm�<u�}ٿ�|�ѿ�\~"����������o%V��՜4���D��X;\�Nݫ�_�����4DK�y�[늩�R\O^�h��ƥ&g]����AbT�@~�i$L������ؤ�p��R��o�f���ڲn��,�\�<��;�����aǄy�8̕�z�F�W���M��B^\	a��1�dQ'�`Ւ\=�%��+ �ܜ�L��!��N�Q۞u����hvR���-�d�*�R�=����s��[;	��g�V뿠��!b��[�z8�(�A�Sd�#4���P��T��Ų6~׶�(�S��7@ی�o_�LTm%�:�v��(�I*��|N�Nj�L!���M]u��(ggg�߿W"\���C��ʙ`b��QH0@�e.E�.�1�ofF��a�V���9?����;r��bCE�탋�\�w�'��=75�"�>Z.o�]mF���o�~__���ͩnl���Kk�ƥ��Ĵ��c��|a�!��]������p��@�_+�T����[@@�8l���X�Yo��*i�z��O'�s�r����|�
eec�@���A��j�C� �p��˅�j6�;dVVV �	����,,���(v"˧r�fffN���H�YZ�F�
��c��N��K�,BN�VF��s�{Da��5��k��}�e-���oH{v�Y��B������i�!cţr��+�%a-�9��-�_��X��o7�6=-]}�X7�$\|�|�v�!b}�����[Y1��!�糰���2��R$KP����������m9uQ���,�����@�!A��C���.K]5���;;��H����ɛ^Ug
���ݍQ��d~���$��edD��iocc��t�^PP@?��`�ͭP��L����ʼ=Ï���0d�cՒ�kkǠ����Y�qx"Ic9|peq�Ӌ@AT�4�>E4�l�
�ifqaz��(=#B�<n��4iI�$�9y9%�i���V���>}/k
:2���./V^�.lm��=<�tm�j��ĥo��YHJQ�+�0��g��_��5U�v=�p�>��Ub�tXH��7��� a�\���6AvN��ن��l~vn������N���j�����|Χ�P
**III@��;��k�;+J�����{f)@�9ZM�"�RI#f��)}e���w4l:�i��p_]{��X�IHX�9�A��f��ꠘ:_nq����2�O�P�n	U���OKf�[�Ѐׄƌ�����%���a~�zF,"���N�V�b%,:��J�����˱��8�#��<$�XGZ�{ t5���F�u]e1���L�_XY��Ϥמ'����p�$�݃��!�d����a�ǩ�}�|��o�l�ş�u}Y'�.f� ��}�2g�6Мt��a��9]*[����R9=�s!�A�.'�m�����a�͂=��EV�d�s
������u��Ug)!(m����xCtր�g��:��x[��ϟT8=��}�x;L���&ۚBA<��a�.�s�mz������\N},���B v�h�>�A����������lR��+**,ǳ�������5 �F+l�������q�I�Ǘ�.%�x��?=&�T�F�4Ts[����L�o�ʉ����Rŏ�N�t\peO}����� Š��v�� մ7���q�z���W��+N] L'^E?i��h�!'�S����e�
pB��<ѱTK(��@0]��aψ^���Q_z�3	�}�NM��{I�M?���#=��yC!��+oW�����'1�;�ݝ-�=|��U���W
rr�*��%Bo�� �=>3n��s~�5���d�lѧ�O|\_^�J�;��9n��"�u-?�T}�J�cSM�Xos&�o����D�\�C�����L�K�_)n�v���fMZ],���Ӿ+i�4�t�Kh��jK�	
3nh)�S��	A}��;S �>GҾ{v�.�_ w{��~ꇼ~D�H6%ăO+|Z�h�$�Vy��^�� 5r�}������Ǐxx�444�Q���pD\�J�O s����*��_ۊ<ϲU*�w/��#Z��G����w��)��h�8�d��.�����ӏ`］��}˧歋����b�'�64�U)H��3Kx-|HC�K���J������@�S�'O���7�ڥ�ܐ�4���1^�=|��܄@�����͟R��Cdxa�����U茚�0L������F����۫YCL�\����TqY	G�7o`��`2���9��ʱddx�p+1)n�U�o�ڗ��U��a�t�2�ak*��bw5�4Ť�GC�'� ���U�5�"��>���3�(}mV��b0���C�1 �?-�>�SF�k;�P�a�DyU�7c~K������|u�,���de4�s+�I��{�XU�׫NdP Kx�{s�lk*�Eqq�,�� JJ��R}�'~�L��I�F�Cx|||ˈW�4�Ԕ��D)F�g����pr{Ÿ�M�X|nn��Y �;� ���9�@��=���֣١�@���jQ��~B��,�3������Yve���'��J`D1ɷ�����V���c@����ҝ�Ǒ��b7H����{sy<��j?pŸ��6�֪�n���x�`01�8C���pW_��*+��ߥNt�B��w��Mz��+�g>ľ�'�s/9�f���O�{�>�J�<�QL<��G������ŗ�eLQ��N�*zx��r���ə�w�[�0��.�Eα�x��O��u��=I/2�Ȅ�AI��H���&Ci��?�:�,�pp�;i�������	6Ұ���@�7��,�;1�2����` �Yy�Ji$*�,�os#�-�}g��U�mi����Jx���/H0�-�Dz�Ő��}.�������!��s{{�S9Gji���h�U��S�0Z_���\�p��1���O���w>8pN���cd����t|o�@�6sQ�����)�M��53M�E������u��d�Q�`K�����r��ôR�\���9&�`>
�D#�� h�\� �3i,�o��0*�2���.�c4��v]5?Ս$��PT
0.������=�L����)�(���aj�(�p�ĤÝ��s�Q����'�ǲ�,%?|@�>���DQ�f����ݛ��IKOς�[���m>ס���XL�[��kR��8�Hc���Y�}����{�ϳ��RVD)����p�Ǟ;<�����va}!ړ�A�8z��(Vyꎣ�I ZQY� �J��b�T��Y�8QPcW�PCGy&`b���t�4a�2�qyK$Nf2M��V�w�/��gW�<Ի�'�Bv��Nuȁ�VA��g�m7=<4$w�Ғڱ����8��M% @�J���u?S��y����7jA2��tXhNg9%]4�a���S�]��*1KKljj��VY!��#�W�CpW%��;B�:s��10���J��z�;��;��v9��P��M�3R���X$!����k#�,66Yۉ�TT��<
i�/ù�VZuZl|�\<�<x��)(\N�ڛ�g�Q�� >٦��R��}��Lu��z�%""���F�q�:P?Z�C��R{������eE�MQjʗO������ֆ���H?�J��@��mI��BpE{	]��;��wT�!e�~VNu
���硖��>�x���#��� Z�_�D$L��5�ez[3��r�Vo�y==�[�i�ޝ�9�$*�A�x�s["�o
�D4�^safl����&���-� �g����(J�a��M©�;1�?RГ��	�]���$!d꿃<�/O����E�@fo�t�/�\>*җ��(pVV�����j�h�ۡ�#*=�v��ѡ@6q6�v6Τ;��gcmX9{�H�xS�'a���E���I�x���t+�e��|@�q-!��S���i�핲0���J����QZ� <͔?5��K#���'$)���� �M{ S�k���w;�L�ǅ���l�E�?�����&GJv8���%<�W�g������?'��ξ�C�\)k �'UUUM���(fjؿA�X�	xi�FWe����Ӌ�)3�%2�F|k�#s1AN'�����t���k�K����z�E��$[�
lVR=۞q�Ď��e��,��m�TJ��a�m���a9�7<;`�3*�g��߄�x�C.)��݄�I�M	rJ68�����_u�G��
P��϶d1�C�/����!�g�>�UlT���m\_�@-=��()9/�q��cs�6���w��A[�DDE���<N�\\\~%xf�x㦡�H�lj���|�ͪ�+�=tx���fSx�� L����>��m��nT� T��B��i���|�����k�������-�e~����֑Tb���1�w=�[���x}�;_F���Q5MS~["�B����諩�@��x�(�A�E��f������Zf��RI� y��֗;��u��m�6mC�� ]��o\��������OQ�_�g��NϏ^��,���~{�9�|$S���Non�}}����7����*,��{{h�%ERRZ	i����	�a@@������f�ff�g����;�@/��{�뎵׾\�-�ƕ�:�$���>�m�;�A�qN{����8�I�w��q�D"������+�o���\h�~��gt��Ӫ��s"��tK����1�yi_8�D�>��x
8�{�;F_'���h���1*��g���a����6W�TJ�O��˄F�[��u�kv�ok���r�� LXL��RQS�.W=�r�v�?�/wP����ߗϟ",Y(>��|6���j�"��nxG4��Ļo�t[��\+�%E��w?dYgC��g��T��]K4��̑k]�3��F4�-ܾ��$�����a���?�"ϭ3�G� � ��������G3�V��^Q7$)��������p<�9��9���iF/����EP�P1��?�+�8f�-;��l�12�/�ll�����,T�c(�����=���R%sB�O�@F�Ƣ$�i�Y-|X$���I�����iN���2�cL��0��\��*&u=�y�2��:{d���I>g���Igo9wX��M�*N%��z���/�$*�_�s�۽��q�a�O=IaT��$D��H��9�Ԃ��=��y;� ���4���ɍ�N��˛���æ�?0���0�5̎g��Ũ=^"�S�y�u�Z�������_��u�|ȼZ��H����r���u�cnܐpe��l����*�Q=��������oH �Vh��I��\�sf���^Kc���9vٱ8���9����w�NG��8�a�����@(�[�9g��f`o|������Pwd�F��,>-��/A�Cu	�<���:�R���G���T�1���{�%������/?q;�������}j��$�\�X��N�"�D��@���U\zzYM �A���hj`k�P2�%j����d�NJA�Z �:��
���Ǒ߂�.��z���tlH�+φ��.���N��1����媞�Vݣ0�ĳK"�ߢnff�5dp���K����ཧ�(Kb
Z�D�4"1�4�xb}�e�w���1^/��:�^+���*���B�����~{�������/?G�]���n����ܰ�~��a
������-�b��KÏÌ�'K$?i����,�-���wԣ�Z� �~�)\#箍������i��J)�)D^���G����Y�5��0y�ڢ�
z���8�
��<����d��������
x��j��k�O /�=,���Ȟk	�9�,�0���aom1	y6�c��ޗtAV�5��q��/�������1�n���,L�_��{�r�)�
�~e�
4�㿊��~��s�N0(+�r�c��������P�������(�M�uuuO�<	XTUW7����eO��^!ϙ�}�6\�@��(������BK;�)]�z����bnFD��~����
���ߴ�\�	._>k(�(CMi���`G�Dv
W��#�wd�S��L�,����L��H�i��&�<�3�в�<IZ���/a��#/��N ː=��@P�#^].��m�~�6�=�%g�32�\br���բ��� N��ʗ�nH�<I���Z�	T�4<+B���e�h��߿��҅����#3�����yt�ck�����z?G�Fp*��뺢�+0n��A���9�<e_�#G>�^��4���������&��H��3 �6q�.�d������Y9�c�g(���{j{"�f��2�j̆��E鰷_�W�̐D�9�"u�f�oV|>�X6��S���s'�t_c^<��p�˂�cq�
�?ov��^�;D�2څBFc���ӭɑ�C�%Y	^o��$�ڲ�4��zX�'%%M�f-����'���JDB(��0,2R�?�*������vQQ 4��˨��-�[k���0� �]�	�i^ۍ�L�WІ�y&Q������p4��epDU<&�o?/��2�?Es�9e[5s\ ڧ*����on��+eo>����ó��7Q%q���U��ow��1���/�T����	w|�<���fř&��lJq��v�X���)Qh24&�+�PB����R�o3,�+�^��Ƕ�҃J�i��P(;;�� P�(ޟh])���x|�117�ce�o�	jy�LЫ��2:�=���
z� ��?��Z�a�����R���D�Z�N�r�B�g�*Z;����aNab�0����a���]b�mζ��Ci�����*#�39�c҆o�;�	1g�\+��Z���@�zǤi��є�v <\�Χ{��|�0�B����^@�$�Ԑ�'_b��~  ��TDs���N����i?�\��xP��4K�6�޹����~@n��ۣ���l�����~��W�c��E&zi��Z̍V��޾|��/d�B�ˋ�����L����'��㙢���Za�S����>��L�g���YLt�A�ߚ7G%��eўS�a�R�oʅ��tUq�q�]�[�w�;dF�m���A�2���?�k����aK�����e�
�,��]?9߽e-n=TY���#?� Jj�0~rW:��6(y9�	1�����9���O�c�ԣQ�����%<]ŁMTr�옚��#��-�Z9�4�t�c�χHC俽��P# ��}N�/�_�j���H9��j��cG����`������dң\*77����=rҬ��X�|2���Y���k�j�n�8+[���j%��ޭ⣹�7�� +Hh3U6�y ����5�Ĉ��S��H}-[y��I=!��I�.��w��3��	G��J˹���7��dR��cV9] ��y�g|P�%w�
��F,�*���$�<����l���+���8�,�x��mYDA5�M������^;�|�}ѝ���@�z�^��ڞ���bwL,q���t�]_��H�^��D��q�ka���mޭj.��%W�9k3�������4>X�s�b�?��ed_n�HW^|���‿�lZ��bf���mu�Oz�d��%�7v�~�8z���������������]���Z�_�-��b�0m��`s�NҖ\�n��V���3��1��t����Y���Z{b1=UT����6���� ��ѝ!/���k�PF��􈢹򰃸��F�|D[$�)t���u�_D�H�=�m\鋱F��#a�N��&y��ZTT�p�.J
�*�	�9_hHH��������M�CCF�^KX,�Bvv��K롉�x��&�G��z�K/�����;������	�y��$�Wg�Z���r�v��T$�wS�]]bXE��nnU�neCbcr�׭iͷ�?S,hd�����%y��`��po����]��{&���୦������XMYeFNB�b��-��
#OT�-Tϧ��k�A�N3��b�3,��~O�g\�QAJ4�)���g��	��V.���@��W���s����>�����ʚ��``���l�t�JХ&k�-,*J��W���A�&נ�bk�5b�=jR���^���8�d��k*_`E���@�
��EK4		�! �e��Rǎ�]X�2��w��vկ��(AV��7��e�E���mBPz��ބ�����/~�_\��}3����\�ޗ;�Y�͛)�mV��k� ��#̰9���������_{����j���JPG�?ݢ?'P��v;����3�H'�v�{;D���U��qfl��\�ڬw���"�\��cWE��.�=��f��ʴ �y�?�H8��Z���MKK�![�E!CX&�Ҹ?�̇����C2��SwwWt<2����r9c[{��p;<���^+��hB1�A�'Ъ�����oQ�*�9ʍ��_���˥��ׇ.;�-��8��E�f���Z�Q�#mQ�4w';����g��Ɲ�vC��~6I!UN�T0��ƴ�j���9O|�>����/Ӆ���"����(�,ҨD����}/���9��
��#���~���BB���~_�z�
�F��3�`��K�!�Gvgg�b<ezs{0��� �<��G���v��ia��|��h!'�_�L�U�?>KHKI�8:>V���	 �7�|�o��fo2y ӂ�}n:]8����3cݺ�gಶ�pK&�b	CǏGW����F�]"�]�4���*�����'1���r4��b��s'/d9͸�x�Jv�B�����ӸC�s������o-�����o��cH4��w��r�j��_ư+��C��n;�b*(K���H�/��T)��c�2�,{c���a��bA�L#q9����a�_��E��a�
,����`nd �C6g.|||�X�D0766�xד���-Σj����-ճ�A�k����ѡi���d�(v���p}�	�V��Pv$N���GU2�,���`����>OQ�[��ߋ ��S)KcR�1�C#���`��~�/��dN� �'T�R`X����٫a��|w05j�<S"��-��
�M��;~�s9&''��bPi)K�or͉�M ��=j-��E�Ic� ���ݒ2��H.)�\$|p@��$����{�F��/q�WU�
�0Q�O����ږLL✔D�
,-l�#��2���Hn�@`w2SL��ښŐm�S�m��DLOqp=����	����	%5acu�6
Ӷ���'Q&�[+�\��1��V888T^M�]1�i�Zl�<�s6���5��KǇ[�/?�;n:�7�>���z��;�Zy�8�B2k�9~�|ooE�e�=-&�� ��/'H0r�+�
D�X�(�9[~H�=T�k��"�1�U������5��a�o��-�&��� M���E�|s��hV��n1Z�E� �Յ�El�����ߐ�y�; [#E��	f�;��А���F�)���B�e�؜��������}�9�GCC����]��Q����0Z�p�J(dv��[�vP>���e��ْ��H�[��)]K�|��ny��F��At����D&K����s�i2����vV�����h?�XO����ٛe�(��?������n�]�fz{q����LmM��Nuqk��.�͔#Ԉ?�ϕ1*C}�sS~��N������Q�Π���b�Q{*55���D���>uL/�F�q������i{W��%^NY��x �M��l0��)((|�,4�I�8T��ţR�	G��߃*C�/���=F=\
U�o����ݹ)Pw��^�υa�0/��_�+b:�|�BMn�ݛ�����F����I�@B���`��4;�G�=��1��Ϭ�eS��)�8��6|�i!�e}��A@��v��NbT���+}����ɋkڎ��>�ʖ�j��eK������o�}� ,$�6�}�#T�j�X�����й���@/7��Yw��w�s�OXD~�ϦJ��.[��wM� ,���I�d�=d�%[$�����tZ*��7�&�NKK�x��������g99��<�3?c z{�Vs�C|g+��#Vq�<�`R�9�O�̾�h�Q�PIL�9����]|�J����Z���U7�xM8䈹?K=���8�b����3v���,�R�̩3�5
rh�&�oVGO��o��z2��T]�D�qxCR��
�g�(_!*�`MEf��ۋY��fL�>B��u~��7��/��
�nO�N���0s��t�E�н�	B�٥72�e�_�K�7:����GvX�}#�y�������+&7���З{�󧾬�+H�jA����ݨ��s���q��Ŧ��T4����q��G�������Cl������5�Un$S�=�� p���U�4F��×�������n���U~xQM���
�|�v�]m�Sf��}���LLr~�Y}Wl��!�*	J��~�_�u=�����I:�b�\]}��$*����(S��`!��S�5��S����%��O���%V]]���c�����s|�)'ey�@+jj~��(�M`���'44���bjj�N����aAA��߿1ii�D���0�H�%���V��$c���f�������S��i�]��7`;.Y/���蹫0Ư!�v��J�u�oyZZe��`b�]�����B� 퉽�ݤ[�I��ӓ=,�ҟ�2}Ų7[�&/�:���x�KW�N!;9�1z��9��n�c��ѭ��~��̓!��Q��bd.�3K�oP��[I&8��_pHf��Y�!��34a<���:��?;��y��xym��.I5�;썿8�
ƙ�Z��:�\�*q�ğ�A���c⚆<�l�����	�_7'�<<��i��e '+Ͽ|�����`�����d�E��5��?ߘ�48ԡQ:$�RĮ���= ��i�7>�;"���r3 ����Xq;n�@ɾOX�r{,_�Ŗj�r�i�.��<�e�o�=��Al�ɳ6���i�����Qae�����~m�K�O�Dn��]������7�@��O� �qm�[Naj���B��s` ڽ��ȈVFV�И����r�v��'�c:��y�Yj^1磗��@��D�*��=��+jLb'�++��Op"�D]Od��ܨ�z�d�=�t7��q���8���	b긞P�RH+ :1T%f����#Dx��x5������!E�jR!%���z�9��AZ�|��H���6�Vܗ�<O{��ƺ�����'Gh��nt�G��AiM���u��y�qk$}e���"3fu�d�UE�����839�⿾��M����S�z����B��k�`��K/��l�J"��677��'��I���e' �Ŕƒ4	��&���V��»DĦ[�݄h$�*�J_MPP+�D"B �z���P�RB�j�qJ�-X,�VM���=�B�b�Z�zV��p�	�w�ؐoN(� �X�BX٭�Њ�9��u8QW)�n��h��6��5����������D�t�\���2�����(�Ї����4 �;�RW�|�V�&dB���ߜ�D�,���;55�U����9���e"O�w�[ yF�{�P;���3������ai�ۏ�O:��B&QJ���V�ow��Vi"��]�7S�����bc�lH��k�lg��gy� �o��+{��M�~~8Z�M��[I�j�m��?%@]h��Lq�}�:���3�4���p>"YK뙳V�iY��Yr>G>�r�md��X��9��m䉣ӈ4!
��C ��ae���qs�yX��[6WDl�)vܳ��¯�r�sԮ�.U>k-����B�}�l�E��k��΀?���(dee5d�p��:��Ȉ���9i���y�qo�G%�1!�$��<�/����j��FZ���zg�ko���X8�/��+���h8�F��I=ٞR���r��"+�Ӷ�=��ys?Ol�������ziB9@��l}?������?]�>,a�%�c��w�L��%�U'*Q������b�����^����wl o�'���o`�D����i��j{�ǝkM39����rᚙ���c䴁�4��)c�q|�9�X8.j��_l}=��%A��������y1	���^R$�	�w_s^?���S�p �ʜء$
6�v	܋���q��[c{��?���ZfO)*b��1}��A;��YE˰V�&��loXޜ�	(��[���'���2��28�4.6�V9� ��ź���J}Z��|��O�£g�a\�e�y\Bs�����$ƌW��~(L���+м�]|N{�X</`P��Jq�,mF��3���+����$��:��L�\��b4q"u椡�I̍����ຮ�6�A<  $!))��������2��<:4J�F}�>��*��Y��+���ˬ�֫�@x��� �wġ�9�:��3�|��P�UgnJ"�4+N��:o��)�ŏ��a�}�x�U�'�BnƾY/ձ��d8묨�FU��V�IɎ�o"1����F�.V����w3�� �),��f��/�;�7�zO���
�E�qB��"'���8fM@)�R/�ρ�{�wSy�ھ/� ]D|w�t.���4i��e�E��1P�����}`�n�Aj���I??aJ*���ߴ���Ŗ����˨�7���{��n��#
�� �}Op_�G�0y�QJ��~S��z�2EgB�Έa5:|D��-�\��"}����)����9�|#/:�Yy����<��%��p4hۂ����v;�C���Ҟ��?ύ��ɰ�W	4�܏/�d6C�O���\��F�,'6 ���r�Z;G{u��,������@��Z�O��:`��N��Z<x7![o����]}�>34��՗�+��ɼ��?������"�P�!�a��=J��I+a<��_��D�����T��1�ի����i|����o��͏��d��{�r$����[��x�m��k.�)����~���n��Y .��-�z2�{�!..^��^8(�݀/��OO[�����5��*j��C��o�u�%?��Pd�����]{��>���搓#:�:q�^
�?�6���}����g�&��-�Gip��2yc떪��U��ެ�$�q԰��l<��� B��;�?L_�]Z���;�G,�:�����ο�[4鄦��(L+\W�hg��6��"����(�d���&ទ�����q��;���0�G�,���4���$sft#�����4��W*|N�/�����]�}�S�1GϲÓ	*o���P@��O��[[�>��:lk����%�?:,x�	��@Ѡλ�`A
a�� �5��%a�������H9�: �-}a��*��Lq�y��ߟ/��
���*a����	24Tea��$�_�n��<W�{��ɡ�^��B6�vŦ�$<�G[d�&�Rp�A&�0����r��1W���qw�B�L�wa4�c�B����.E{Svm��>nzJ|������1� ����>v�בfW�ܖ;|*�l ƹ�ak��JVq�����G������+�leC������{^_-���8|y���"��[n V��+Ӎ�ؿ���"����>u~�N��+|
�!bsns8�����ݥ��������������l���,*�D�X���־oQ���wMm�i��J%�qK��N_���(����z�h���ys:,h�x?*�S8{�*�G�P�����h�<@�N����Nk�k0߽W��׹��ZqvU�qB�e�?ێ�ޅ��� n������5��	�~������AP��u�m��B:�2ǺJ�/�|�Lguq�T�Л�縐����� ��5��A0�w��%(	v���"��|B��"I	�b��&\�ݥ�����G��+A��#����PeH��)c4m����!��'i4��om&b��s�T��G:!�kd�<�Qs�aƸA9���xu��Gin�rZк՟��G��$9fk��<ԑ��0~�����0�ƙ^��6��*i%���e\&{��6n����}��S��|��C!cZK��l8 II�
����J(��V�qd�R<�d��G������k{m�׾֤Q��?�E������F��u3��Dp��a�@s�H���n/�$d̮�]��w���1XK+��{Ό�Gx���<�P��,m%�	-�RFt�tlp�I#|uy��!���T���i�k7]��L�Dm��^��:����4O�7P����⻹&1�4��Z�|�W?����}�4ľ��ް�q��B����W�M���.G%�\�h�g�����q�z��6�+�b۩L�K�P<������oI*a���5Z/�10#	��%������e��ٸ��V����O��`��t���]���e�b^J�H�w,m�mR��^���M���$U��� �t�+��[�2���a*�xT�������h�%@�ө��qM�냛0�r�W�Z�*b3��';���{�$���	�C[������H�T�řd6}���KW�~°�7���fuq'V���&�;�i{�n�LC�@��qx�#��HV���͹�}��_�T�;��(��զ��� ^�߿Uw��DV����g;��m��=��{���4s�Ai4P��Vη�[�������{���i��ߛ�
�d��F�:��,��D%n�6Wכ�{^��s��ȅ��G ���7�M��Yh�����;�؛��B�|ڱ�gd/��yn&ߎ�ܴ�G��Y�j�����پ���0:jy�P�톒�Q[F�����0�"O�,0KCR"�
&W��1'�=�/������ʝ17K���J����Gj�Q�%��^����1Y+'jC�D��$��wA��;�6�cnnF�D�%G��x�/&���<l��x�}�{�7U��s�Wn���GIr`�uF�C�=�}8bR�F����f�7.{�e���D�e��F�[GYE�?��]d����	��<~b���A�L}�C����D	\$*��������M��{�gmik���z�>v�c-/��U����? ��rt?�TH���*���.܎�?��f��ޖ�Y�Nbsx߇��;(^����s<��Ytl{؄��6�z�We-�2�?50�� z�*�e+��It�w��[�#�������j4�rm7�7���݅�ݿ�:]�*��t_O{�e�����}zQx7K?��.GDL���5���iP�s|,]�:栨��+�d�4?�z�~�ؒ%%1xm�tN��S#��7��qul����l�6�æ�;���!���ʙ<cʯ>b�^�u�����xy{W��M�HK����d����Ez�����]��
٣�8<�,Ȗ�"2J����^>|)A>�0�`�,#�R�v�_7��j���	Rw��g�\���F��ן+�uo���
�V��ti@�W��E�'#�G��7Aa��PӫN�G��练���%��Vw�A�K�A���i���J���H������m� �"M�%L����Z���>L��klB�P���)�Ɇ�����Esu�*޻ӈ>�����f�'j�w��,躺B����%�%'��D���(�^�'r��c��@v�(�T�Ԉ=�v��XS�=��ڕ����˸	�nRB	8,�ڎk���/�y�F)<K����y#n�lt�XYi�9���_�E��NV�䜢������͏܉�����.n.�!�g;��gA�����>�)j��F
��ɭL�u3�..���pgJߋ���+�cs� @&�n�Q6oT� �"��me�n���-pJYx��!��u��C�5~_�1��I~��������j���h؟:�����Y��|	����Z��N�= W���.,��/�ɨjg�Zs��d���Z�;u[��#t���J�ó��
lka��'��������y�S���.�����cQ�MV.�Z�111J��n��{�o��5�;�|������e�#�f5LozK�茮/	8��|g�\����Ĩ9�Z�N�ʆ�Uq�5�X��tkn<�7�R��j&���]�������c1-#�#>L9.N�-��/*������ O���zMß����fڬ��ڜ��ښ��2�h�����6G����m����c'��a���B��c���=�5���V�zN;��Z7*���)��"ܴ8�yRޜ��v$��t��t�gCs����a,�;�,L����:7��#�+�.�V@��z�Ѹ_;�谌����qvt� N�	y��Ӄ��z# LH���͗�]��q������,���}t����"b��!�k�+�ut>��[�4�me��E,+l�,G#	���K��IAN�7�w2�wH��~�p?�W�-r��%�\�ϖn�N�

�{��!�X�ՠ�� ߭��#/Ӳ��$w���EN4�y��g[���,umJ�ܝ�O�Z�u���G�$�y21��LmSIh�Z+d��?��wɤ��<���OF�F�s��^���1�������7��� � ��Bw�Y�����]�ڮ��e30�b�"�T��x���Hy���M�}�ߖ6�I]�b)�o9�������h${�9���	�E�ޖ��@�Tۭ�B'�%��/q����N;H�"��NQy��`[�����tm��m��?jYi�s10�i��D^4�UR��p�+5%��RӺ>�٩��}5M{P����t���O����/�k�3�U8(UU����s}"�V���E������-V��,�y	��v�L��qͷ.�^_�zmO'"��{o0@D�]|aB��G�I�jBЫ��A�'W��V��I�ecV-qBח)ƹ��w�2�q��v��}��v���Z���ֵ<����)ϵV��"���5&�"���P^�3YI�b��ܪ���G��~�����B��I����p��ҍ׼L�Q#���#�[S���:�����RU�N�!���
V�PO��n�V;�����~�5�� �X���'"�<!ť�ٗ��Z�+�7h� 4]%%G9�볒/������m��b20�qA0�,��ؚ�����==�$���⡜�&���2�uy�L�	�����R�Ǻ�TTi+�C����;/�*/y=-�����sm�3�NE�bu��FM�������CC��͎�6�98u)�^�����5�M��ےS�P�T�ZU���o���a��AJ�1Wj�C�{?��l5=��:;�}v�^L�XTx�l�P|M��DLb�<������H��?<��g���E;a�|h�a��t#�T�����[H��٘�� *{B�x�Fv�ŭW�ӿ���l)Г�kl5F�韄M�/'�9]�AR_ u�o���
�yRO����ױ��U���V%�8��(�ZV'�+�y�U����&6��v��R�]	4}U6E�ξ��z���Z����]�BFN��S�a�?;���˴%LNn4Owh�u���x��>[~[3���7T��������WIE�(u��@����Ϛ[3��n��+��	�_�{��,�lS��.R��#�m[��N�C�-�աZ��CUy��Wf���;�5��K��H��`�&���k����.�؆G�6 >  {�$���D�f�a���@E�Ɋ��	9�eDئ
U��cx쫙����H?K�6A�����=u��f�%�e�B� �ۼo����h�?�ɵn��4�eF��4[~HJ��<�����d�=�k����+��	�^!���}��F��s��<d�!t"��5��|t�Y��U��[��(V��tn9��'=S}���q�����>�3�0�!��n����[��p슷S�[���.Dg�S��!R*��%�V�QtRj�Dn��B�R(@ "<�1��~��ZBV�)����h����|΍�l�������=����x��ݎ�a�=�©~�� � �`s���vA�ۯ�7{FP�h�A�����E�_���<�c�<�O4���B��U�5�L�Y">�#�H9l=A E��@�t�Z!!!�X(Cxxx������e��XAB{����\����b��0��B,�b*!:;D#����<"m�����E�ʐ�q_�w3jn��s83�&ټ�A\�'��Pa:�ej`K��ے ��k������"�z�;��+�,�o�[�g���Ǭ�h�f����'kز�䒽w��OGA4�{�$2ۇ��!�m?�x;24nOQ[�w�R�٠BiQY���h3���\%�;fRKh����XU�C\�OKw_~������������3����#,?�>v?�
*�j7~������cK�F��ޒ�o���+'�\�޳�ިخ�p�AE1�����)�Dj ��e�s�"f���*(�4N]���'�}U�5bߗ� �M��x��YJū���z�:��1��E>�o��*� ��u��V�<q���eB��ǯG��&η3
��f��F����( �W�mvޞ`�_�eq���FPfE�o��mb��?�D�p�2 �����^111��N�b����]
7$�I��2�	]����wp��&��w�����o���A�Wj�͵�&^b��F����`kWGV'$g ���0�w��K�@�bZ6
�2��&F���X!g84?�n|y���A당w[����[I�� 3F��#<)��:J"���7'V�̪"��<�i����(����Ai�+���=��������2 �?���ZP��{h���h��Z���S�e+�p��L��5���,	�M�ܻ�NG=��e"_�U����c*vbi���8Q|���1`�9|6YQ@:��Ɲ[��'��JD-��Af?1�ş��6=����O����9�N�#��!��[SS����2���|�jW�BӜ	�����Ww��voa+H����>�,LL���.ˌ
j�@��ݜx�O���(F�Xr��w����U�LB�}�D�_E%
�2��i:� ���:k�����R�3�Q	0�\�'F�J�듀���2���^�mX�L6EX��p�	�D��8��o���)��F��lH�t�H|�!( �q%�����	|mk=��/���8J��k�Vд���vf-���� C�ش�?�9��O��� ���xn�ܲ�0�-��@����]��z��:��WRV���4Z�
��IR�W		e��	��(�r8���fd<��r�g��r+�P�ϥs��CC�9)�X��N��R����r�o"S?0�#T#uO���AƹW�ߞ_��C6?k��g��]����0���!���bJr(�IZ������,�{��1����(�q�8���	��<>tM��e�5�\vtǣ?9�QA����+n+mR\_�#�(u.�K��2V�
��.UE~�@���o.�^8�;��mPb[���ﺝ��o�UB�~b8Opss���O��[h�P����V 6�n�E����.X�	ӣ�e0���	R��U��X �t$���3" �����}����k���y�m��̖�U�	�wEH%��A���j�D�![}�[��QyA)�x=��<S�Ɠ���84n�o@���E�уޙuMM����B�e�T4��V��<�Z
��׻[{)
�ݣ$��zs�9�v�&�1�%-�y@ψ�����W(��l�q�O�>������=?r!� ����@�|2�V���SF����0<Z+�J�.#��3�eEfy�)�@ �����zɈ�z�Ԩ�+���_�V;�c��)%��i�A�%6��;�[��E�<|m��r��,U�6�v���!Eּ.��w&m�sI���R�g
��jCa��dU����ζ����ɥ�("�E��� �v�m��f�7�����LG���r/GNzb�w��c�?FJ������L�p�����·�%G�1������s}d;�e.�8.�cx
ysj�5��T���m��XOe�]-ذy��иrLJ�xmǁ@֯��LFӅ(<�^fb�����B��c[s՟e chc��l����4+�о���^�P��9EvF����ɞґɾ	yn�u*�y_�5�����(���%`N�f��vzSq#@�l�����)j�7�����s�������q7߸�c)0͓rב
�B�Ps|�2ۑ�؂eH}U4�Z�$�ۘ���Fg�8��3���F�"g)>&�H��r�gub�"�&��|F^3����?0P � ޷�%��I`L�;�ds Ͼ�g���w���F�!�о���IȥP����81i!��ļ��d
~���WY:&��O�١�&�N;�E���I��8p,@��w@
��|��g��}�H�v;�	��t��r

�p�cxR�Z1gMctkI�X�m&�K��2�0�L���[����k����F�WӡH��f���g�\ �X�x�W�c޳�yc�K0�[Z��\J�π��g��!R�J�X�]`���Y�Q"6��.��3�*Gx���JGQ�y�@q^�H����Q�TPǕ�� ����NH�n��ڢő���Ik����n��9�oh� ��:2�Mp��������\����@�|w��0K���T��M��eo�q�LX��o��-	t�J}��'�u���$�x���k���z��_�|�j����Dq_��;��]��r/�:�&���b��7��d`|��n�{�s��X�~P
�����Rpم����}��`%�];JVғ�x�e9b�����>��;��!ϝ��#g�(�͏N�
4�����ӟ�&��H��N�������.�md��J�!R�._�&�bY��6��c��Kk�����
h݌�����.
��ABoffF������C���&��}}�˱ I9������i���!v�����w�lY7~�JB��Vxw$l׌��>�f����bd�����"gےFH���>*�	ú�ٹ�S��@0WF	''E��G���`m�)+{Kf�&������}o��͒�V �Jml@�O��h	\�ܒ��$$��K�j����x%mm
O��y�9�-_�+�ȑ��x��<k��P��.O����`P��Cr��s�M�
���@�0���P�,��[V{f0ۗ�*#�0+����]q��$%烀�����c�[&&<P@�̡�%R���T�b�V�K��FPO���wnVW���ul�ʿ`=��e���w���0�;��<�^��&t�-ӈ�;��-�ϓ����C�F�z�n�/M�M5>d��; 'IY
]��3�]�r�E�_W��MK�	�-�ڌB�#:��%4��7@��ғ�ۑz����M�b"�:gi虑����R��� ��''�L�QU\c�|���'p��z����)���ޛ�C�F�Jq�=[��%$BY�	I�d͐�Ʈ�U7e�"�"dϾo���}����2�s}F���z�~�����}W��u��,��>�\cB�Uf}�W��'?�j%�C`\P?��)8�ysΤ�]$4�5�&�͵�S9}��@��P�Gz�.���j4�H���/��<"|c<bB�s���Q,�	��eW�m��F9�)@>��. �pT|�\��C�3ͺ����QQ���NK�_�kw�l��G�e^OٔC��8ޏ' B}9�8\y|��bׇ�T��;�Za��8mn�jy�Y�=8�{X�Z�gM����Z|�����F�Cُ��<�(B*+������|�aoo����6�{���Ԉ\�ζ�6}EEE�j��U)����A�.�ԟ��v��ǜ�7�d<���&����&�'�mq�ˮ�:�170S/�Y�>�>hI��-Ӽ�3WX��i<�W<,'�ʑr���iŪ��d��9z�r�\,C�����
�s�(������8[ޕgETI���<���]T�J�-�O�Blq.��v�s�u��9��J�:�ˣ�&d�����H��w+$~���n�<�l�aK�"�C�ۥ.�&��6�Wg��T��r3L�<��μ�e*odk��_�/�̵�ڃ7�����`��74����Ӽ����I��Ĵ�5	��kٖ��]*esunl��%]E�����?<�zz��y�'��<.~z������ғ��i�֏wA%���)yQ4�ᅡɹ�)V�6!�/I���wغ\詧� k�Ⱦ{�����}�Tv~p#~��#��R�R��R��Ւ��[O�(G�	,�赆�_�<�K[��1�\ٵ�����{=@��A���
0������K���\侎P���i��ȭl�r�/kϰ�j�TF��9�EM���'J�M-�`�l���Ǐc�
�yTTd����G���%\�a`d�k�"ЍN ��l{��d@/E�x*T�9������[0�}��[i1X��$�FZ;y���X,4i��C#	2ۋ/�O�	?k�����{v�ض�Yk�)�ޞ&Pt��y�z���C����h�j��I�8��Ç߿{�s8`�TT�#�mU'*����޽S�GE�1�����j[�?i~�q�]��
���0G��"��☎)��z���������2//�{iޤ��8����K�>������utt�ߪ�LV�]����Ҫ.;�O���	�5�?RW��B�0X��qu��R�{H��b��,��ݮ�9L�4R�ɓ'{���$��rZth��*\@+!=�D�%���x���à��ܢ+ҫ�Z�JH8�o������)T}0W��Wm��<N���hA�]@����� ����f�r	�/��%.����֜Ls���<�/�*��M�{�XB�̝"(a�y�xt���*��j钟�Z ����O�!�c7���05q����ׁ����������f�|L<wHӓ�I�2�Y�Oii)�> %T��	B��}IM��t�#�Q+�p*���1��O�H�kK�?O{p��eW W���+��%��U`[v�$���FFF>v��<��::(4k���͏��sN)�Pop6��Mo�s`ʝU��]����w��;�o֛�q��~�v�� 6I&P)׌������_y̷2�O���k$��/s��5��	����es�N�?߿�yZ�j����'7��ݗ0 �֮�p%oo	�n,�1�<k~{��#=qj-�B!�\n��.	���w5�x��&-�
��{V�$��g�Q��^�L���Wn��n&T�r�&jƭ1�O�y�~�
,×�W�Vd���.�g<�I���`ll<;T&���A,h�3�~'4�y"V�*��U񽠿�L�~�&�S"�͑��f��=�{��ba׵دX�Z݁�0�^�d�[������UTT��i�+liYY�5>�G1! �Q�"$yg�
�� ۗb��f�O�t-���Xt��Vˡ���4�-���{3���_��B�s��tjt)�H���H���<X���a/s$ u�}LMK�ew�{1�:9;{�N�[��A���U��?�������������f=�e?�z{�\W��ۤ��i=�x�q��ìbm�m��S�a�����qKm�m�4���&t��.�)b,�����)�˻6Z�T�-n,�����r�㐽F�R�b�� �]���/�t�/\M��hۣ�zqq��nen>��S�s�rt��%�P$�� !ψ��"�Y�=�l LXXY�wM/�Z}8Fs����+�H���N���Ѷ��jdiG��_�_�����ִYO������2�4����+_��J�s+���Y ���+E^���m��շ6;�w�'*+����tߛb�nrZj��M�� 8�S��N����X�D���b ����9��^ԭ���Y��b��c���	?�)��:�����_�~���jF�Y��\�H	�t|ⳃ�P��p������:b���9��D����� ���UVs��{Ň����ֈ�����d��+>U�3�js������ ����OZ�u�s�SS�,3���VBR��y߱"��C Hg���<�{/��h��¦]�O����ɔp#9�ʢq��mR\�����w��B��D��i()K=��<�e}�O���-���:Rk�]����t�U���>x�,�8�0Ֆ�FȚ�+f������O���Y~D\]��%��m�		$����(B��VX�2���B�;pO(�KMU���Dl-�>���״p��y�������&｜�|��!̵i�(�7˚��g��	�M^N��4�`�� Q����P����>8uafYn��G����f�>|�F����FM�������d�/��/(��߅f�_��%�xke��z����B=bi�]�z��1a�� ��iV�1	����#lt�� ekoKk�d�
ޛ�u]�]l~,G��Ս��*7�F��y|�(�R��5t�yؑ�9����м�9aI���a�u:Pv7�'9@X��gs�^����� ���ܫ����oC��e��t���0~j�W�1���^M�v���Wm�c��|�"*�}��쯇ܡ�7f��utt�N
��p������恻g���xM���q���]�ڡ��q�����ef
�y�c��?>�X�p@�ݙ�������q�kX�v�>����$h�����8� ��|����ˠs���WFc�r����Z(�0�q.0j
�tE�:oo<H_���
I@ej}�8��M���<�kG ?�i]~:����ԇR��Ο]~���b���@;�E&��|�Z�%<�G��#T��`-�� ��ZE�K�b%�G�]{��\js6�x��a�yF������SRx���9�EN˸H�!�WGvO� �'��\1��2��=� �p�̺�,wsG��j��X(��ģ����{��⼤�_G��dK
BV�Y��Y�AaW���� 'D���w`� V@8�n�I��?*��� ����: �c����RS�(:--m��-���IM9VÕ�/ o��@�PN�yAH�$� �ǻ����울��g>�>Ǫ�!J �T6b��ۉ6�%??7����j&''룊����PBB�GS�#�ܭ�j�%��tw��cʯFEE劭Ex�����f��� ��O͏~#����*V1����{ɠ��u�|���?�ʡW�'�7z��d��.\�+��~IM�NϖC"�rL��l|ρ�� p((d<)� 4��&��L�'S��:�?��R��x�uxM�j�J�'݃�Y�E�lu���zH^��/*��"Tͯ�h�����(R�yH��n�C5�I�#l��6z�:����$���A|�����%�2x>蚤$�_�D�����4�]}U N��{v�$'�����֌^[��E���x��tE�̡vcy&/h7z.YC���|�P�lC��	�� ��ki�<ݍ�X�����w,��ʉr��=Z=B#p�����b ���	�_ �����]�a_Pv�v$)�g�rn�@%���t�Ü4��D��{�e�l�b|cU�ڷn�G�8-����� ��h*@�4��b�.F@�$����VA�TW��Cݓ�?�#���/L�|���%R;=T~ ��P��H��>�����i׎�ʒ
zu}���jg����Su�Rvkkk_��8�fܮ��j�� V����-���!z�P
�#��5ݒ��gA">X��E�e��8>��KG�OOOG�����
�jn �|r��bn�$���?W �0����ޕ�vvY��̻�'��~��￱�O� X�A�#��ș��K:Z6G]�)���zf�w`7��9��(�`軠��]!'`w=�}��`��=���\G��O��ʩ�#T����֙����g'����8��7k�����'�c�7��A�ŸV�k�zo��xB�/�yy�,�'�㏯c��[^��k?T^�K���d�,�l�\�[v��}��9;��g�?E*\�hC;�xru�9&ҹ�Y:{4ll]�rJ�Ն�UW�������d>��?2������x�I�g1\V����^��_rDݯ+691�f�W}����fm�B`���a�z��;�����e@����l�@t��؄�l���y�~�Yh
�͟���T�jf��b�[i>���#~�i���khS����z?~�q��G����3�F<�[XLȐ��ؐ7�H����kLL�K̞:Ay�� �=}/�|��>GCљa|B���Ԃ�
i2n��RM���QX�~DϨ-.�"���:]'f�������|ߝު���y��0[I�n��e���t7��$�5�]��y�E����44O��jU�t����Y����y��v̕Ӕ�(I���%[_ֻXR�����q��G�E����#͂����@��p��ln�mKbG��J����>/�%ޅ�mR6�MO����
Ǳ�[�7N�o�m������D�՛#G��v�;�;4Hf��5T�|��%�Y��R�Z�36�����q:ݧ�z����Ufm�g)����K�����Φ��]b�iM��K�	��M^A-���_ۆ*�޶%p�-|%�s,�TT �c�d��0����RVOQ���/�E!��U���:2��g��6�X�jap��p���ӷwvQ���y1+�t8���M��;�����3L�ޖ�O��?Z��� Xs�p���t��bWS���r'���]m{+$U�(k�aTʣ�V-u������gWW�)�6<VLMU-�@M�A&Kx� >��is+^����{�>��v1�X�e���C��r��wmڞU�\����։}��A��|��]��*x�t�*vL��e �*Q+4�a��Y8�ms������Ĺ�����'�Wio�~L�I�c�
��j��9��.�\f���'�D�[�a���j��2��N�I4�(�2��6�993H�.JU/,Y��^ɴ��cť�_���[_�?,�چ�����R�W='َ�ța�bLɢ�2A�uR���o���~-��7��	��di�'U�#���!�0���P�[�����Ǥ��=�:���g�M�q�Z���M��g#�\1��Ė0���1ܺ0��F��
F��?�e1��])	Q��)�^}m��:��7�qrRwD/�k��0��+�^�9n;��E�,dC�,A�6>��ܿ7��!�g��z�~�L��ucsG��L��u�|k�$�hm,�Q�A�viE�10�v]m� ��Q�_��,�s>���(�}�H����מꬦ�cq�Z�' ���L{0��>��ApS~:}���
��G�����G��ͳ6ح����#h�ۇ��^�vl|PWh�?�'�+E�l����v/�#؄>��D�3�
*����+�u:�*RU���ȼehZq��E���G�Y��aQ6Ʊ���{lB���x�/��i"r!��ǎ|���h.��r���ǿ~F�~ƶ���~F�?	7)ߚܐ041R2F����1R�VIS݌�tKd.��*ۯ�M�WP��BAyu�����*�$����$��l~��-K��X��54��H�H�,$�#V G��n�k�	�2�K��P6��a+̸ �0������r��M�"�n��$Zb��6/���m1�'�V�`##���]/Q�u�$y��������m��A٪����&,�wZ�VѠP�`�U���hl&�ekЀ;U|O_��m<�L{3��-��7��@�T3\���y0��(�_��3\߁�tG�~�~kB����@�r�[����3����A�Y�5�� �
)[0��Ď}�(x� 8.!O+��x�d������Y�@@���E�����,.�C�X���	q�B.����w o�4�Ln\�c9��kE�1#-���7�^KO�~������?xQx��U~{�|��xV�Z�T�i/����� gqHZܸ�P�e?GM�\��t'�k^`��Tfa��{��J��Jn2n���*U���s����K�{����_���O>�v�Bj#4��G<��d���ȹ0��=��������:�/�S#˿[�v��{ t`
@��� ���!�+��.+���p���"���.�p &{guO�|r.�E6���5�1�q@� SʹXa2/��s�[t���~k�Z?�W�Ub���Ucǫ���qy]��a�_|����7h�_Gf'p�d\[��_�*��p��h�C�_㘋}��ٞ�d���H}�݅�`�/*
�<C��+*�90�O\�jRKR�������e<�%��4I ͔� �s~����o'9�#�jl_D����1��vt7��<h�(s|_���{�� Z�ɀ�x�oϊܰ�姓��}��Rq�<j��?\�e���,�������Ղ7_�v��'f遖��C�0���~�=7�*�g\���cr9��#>�qG�VqE�����<z�q� :>�0�֭D��t\qkPn�fr�Գ�i"��a8�	@�=���6hG~Wq�7F!A:���'�$����������-��4i#+��0,�J�$�+�"���R�����v.Fo��=�T��O�b�6T�ܰe8�����E+�TB*��8tB��Ł���j���嵕�}-+�eA�>]/r/�®�I�fahw��	U.�\��&+�\�n�l��|U�L�<9��p�#��_h&I�<
}nOmEr{�?�*�a�0���-�4ް|��*ݑf�Cy%|�
�ʜ$n�����E4���
���?�TG;uP-͋4�VJ�Z�ڵU��x��Y0�}=�"��+��:�����r\nķ���A��ʸ�F�!q��w�jcs�
c�%�̵b�����c�Ǹ?te`�5�B?\��[��d�v�l�I���ꂎ���E�Ê�L$��V_ ���򊢂��E���vk3qH��W��S�%c}�&���Ns�J���
�9c�����g�`@V �jvK�k}���a�t7�ޘ%&j���@L��_�]����C�{ai��������՚����a�V_&�^���:���co��Dd���zhh��[��~�a������h��&���T� �
�+�ߘ,�|d.ҷu��hNn����S��ЎƼ�L�.���s?�[\��j��q�#���.��]�����K�7����»�˔�s� P�w܏j/�Y?P�&�����t>�>�Ђu��g��u�s?���\Pu��(�w%F���C�n��>m��t1Ԫ6�w覀��\]�:K}x����
{ՇaFל���u��>�*m�P��I�V�R7����:��r��eç`O�Ќ� B{J>W���i?��T;�o����ܢ�t����
���T�W_݇�B�� �ӊ�]�$bm�<�?��_a+]��=t���k�W�:
em�B�����
�i��Y�������uL�m!��9u^;�5Ī��*��+�!eO��A�:H����:�{��~ҳ�4�~]X[�P��7i� �W&�wy1�.�0;��Z��66oY��q�h�7~;�c��!�|@S��;�ҿ�6C}}�M�P�}Q]j�*����ks�K�E��P-`/����1�X��WX����Zc-p�Z@���_\��h=����/ڧ��f��=���(H��|�`]lŷ�����)�\o��:�jU.6�}���O�"Y�����*��6��xO,���fN�%��p+�aw��}��1�ˮnD�iEr1Ѻ"�Y�NZ�QD�ĕ�+���o\�R����4�T�¹Y+W>��F���,�2Qh�X�@ASO��g�f80���o�}c9}�.��@g?a̞��GY��.���H
3�C*�&���]b��ػ�P���{�қ�#���di�����ڔ�Qs�-G~��m�nb��϶#(B���Q�ޔީ�KC��G����'e�M�?�,�E��2~"��K$�z��� ���X��x��SՆ�M���}����,I���ܞS��%��nu���-bHzO]�|��xE�`Z��ܫ��:}mgG$��@�e���|���k$ٻS��?O͉�#������.�.r\�������rڷ?��ZT�}ycm���mg�'f<��W�}�I.�j�e����w#�����z���4^u�+5'مc��Rט����xSE�����×T-t�AEE�5W�D%�9�rD3�d9�k�z�A���_�z�E��Z\<�P�c��>߱��\�l�2�ة;c_�dى+�h���U�b"N�B's�ҀM ��.�|�	�W�t�b�!@��5P��U+��-�Ht�|�#���Ⱦ*�&b�=ѵ0��s����jn���c��v㥫��C+�zg��7���io��v4˷��G���ºB��Z�ϕ�ʡ����q� P@����B���@���{^jH����	���US��	yG�Y	R�gp3�G(YLy�vN��_�İv	��v�~�L5-ՓofUO�J2�Z��
%���|;�NTTK����Є*(�z���|WJ\���ϧgZ%�~��䧊f����9���m�M��T]�\t/(啫{uj��N�{vl4�^ܜ����¬ё6E�G�%�f�6����s�aL�5�w~-E��d�f���-%�#_E��"9��AE1}�r���%PVA�7�ܦ�&��#�:3��y��Έ��F���C����?_Q��a���`O�ț��u}2k��:g���m��nﯤ��m��@`_n������3���*钫��Ub83XU	L����n9p��Z���ɃL*N�������O����r"w�,M����@��������"R�ۣ&n ��Q�n/n鹌��$ȣ�¹�F��u����s���=�,*����X*9+���{�\��+}��4I����e�c���xgX ��d��[����9����~����x���g}��T�gN!�̄:|��������v�e�;�+��j�����a������L:��=�Ϻ����~R��E?PlD8�t�œ��s�<S��q�^,�wd�0�;��o<������j�W"̨m�.Zqm��}���v���Z]�Ʉ�{�� 9�Ϝ�};���ZX�}�zď�S^�%���q��K�H%)�_X�e[8���еc�3���Q!^'vuL��}�بmh@�'�TbB>��L
���+�\�ʅE��m�z�3�����_o���,>t�؋W�Fadt�Cljia�[�+S��3ןL����,ۑXtc��I�bZ(Q6�� �}Oq#4/�f_͟5��z���0νK	������zXh���h�e�EĦ
G�p� �!�&�w\[x7���~_Z��G�'n�k�e��m���
�җe�IW"gz����čF�	�}+`�����^[���md~��6������LrD����RVu�.J�)�Ùe�	�9�]�/ݐ;w�X#�Lh���O�R4��жʗs�#�qJ�m����+nv*�K!ծ	t����'�g������8k�_���o�p��7xC]K��H��w�~��+��^Z�t��U-�w�ߨ�t��i s���[q�ᆎB��1����<�����{ɶ����Nq����^�� �E�}�P��r�2����a01UTf�GVU�QP�}�����2�3�a_	�E�U�B����k�;h���;��|�}�7!��ь�K�'�l��8���5���������7/feW�A�t`~�򴠡@�̹=K���+������p힚e�ԙ�|4o��I/MM�Hk�Kȳ��ޜ{t�9���]_���j߻���xz������
;����� 萍n� GST�9;7]�� z��d��+ō�m7�0�s�m=ăؤp��s%�.X+ϲM�_+y�C���Qq�R�ji������נ��l�~ՇA�Ů��EK^�J����[�"K/����ۏw�'yB|5�~���N��\bްT[8��k0�E��V����~�����F�^7������'*��K[�ɱl��L*��Ɲ9���o0}1JA
�ԉb�.����Y���Rϑ]��I/�M�|�õ�i	��[f��v�N ֈ��{�LNsx�
�E�0��kKp6��3^R��3u�K(P�)�� תװ��s�ݻj}���)��z0�4S���"c�e�����=�fZ��iA=�GcX����X��<���go���rZ�C�h���|���ԋ2�Y��#c�2�E���\��>$,!N��;}����׉�41�kh���ç�*�$d
����N*	���몷��F�fU���vr��<.����H�^7�c2_�p���s���ŀ(�	�x�}�á���=�d6 ����&��%�?w�r��;e3%뢪,�S������΃��|���J�E���ℓt�)��,��^6����̪t/������K�W�/�uݚ�6���	w���S�Z�P��9�R�ܜη��|kK�E���=,*t |fg�[\p�f�$Ο�E�,"a�2�\�^�ve?<QT�&�z�rE��b��s�d\GЊ�Y���"΢���!��֞���W��!�z�r>t�&���v����h��f�u�\��<��%WƱ�Z�Y����,�7 ��c��J�K��l���u�˻�h>���?��xV������L�6	M�(�"�g���2C<$�A�9�>���_m0/[ra>����{��x{�Q�s�k8���|������~03땈���{=%P_����$SX�2Ӫ�G4��8��*>
��)��v`Ik��uu�_�y�׽�p�����h=
+?de�+ܠ���9��}n��Č[�hR��㗤�<!w�կ��D���*Z�^�V��O�З�N
���.~��"C�oBZ�׮����>'r�F�*o�Ԝ�V�������P�� �[o��^���w)=
�]�@F�_�4l�>�)�U�6 ���� �pO�X����}��R�`�����m�PJN�\��.��1\���С7#]'"�5�zqHX ��q�w���*���<z�ܖ,ǋ�Y�▾Mw�N$�]3������)�6��~�~[�t�����	Y����X(�m�7
S�����xKO�7r�����S�:�-��xd�>iϢc���S�e�r(��T��o�7P@��Fk��Q���'�<�D�}V���"�W_�V�m&����(b�;��e�P�x�֫���/7�bUk��n��.;-f�v�<�z3SM:"�n��]g���g�����T�N����T��o�ʻ�y)���W=�����f�ʵ�!�4r�7�EhS�5W�}�xݬ:4���T�N��}�U�5��#M�eA�zf���Q�=:G\&�O�D�����o��n�-*i@-�?������g��+-�&�C����8��O���d�[�<���T�U����_ �4�3?)���X��y%��@���ɵXmQџ�q�KJ�pfU}��OQ=J���&7@E��^���-x��ٟ��}'��:�a��C�
3k�Cn�1�w� �,��k��i?G�G�;s���?Îa��z~O�W���H{#����k���ʔ\�H��׵W}�S5�SL�*�v^�!�-&�����/6�eE���,O�2�$c�y�z�T唎�vv;����1�>\Rp�q�����T�%(A-�.]��g�4f���v�R��S���J$�����S��R
�Rט�ʟ���h�U�U��p�ma�-�G�:�&G��,P�8-��C36����s�/�C�:i��(�
���fdΕ��.�^���ߑ��@9��|���x�=1�����O�H����bm�MK�͸���_8��ӯ���d�+.o����	���7_D
\T���4mYw�v�X�b(�dK����&e���l���[g<\�w�A�jc���\zd���o���$~�z`���1����G��ns����:�}"M*m��ߵxW��	������LP�R%Y�P���-�$�z����w�WH���9i(��A�N��BH�
�����%���C�Z�'C��r(�*4g�� ��#�ְ5���(W>�>�s;os}ڃ#�nhIUdKע������&�L�t+���WT��>B�taƅea-�i�����.�Ƭ���ב\����^qY{��^���jN���}��1�x�JI28���ޓC�ŕ����}G�s�,�ܥJ*��,Y��n��/\{�V�֤p���!
�HLL������t�]���f�;c��n<!wȊ�*�ґ����R�CM�\7�����ⷍ���/Jn�L�_N��^1�a��i=P%�=WW������� Fr����lc��sSR�^)�K���f/^E�� �&�H�Ȉ7Z��G�Eo�a{l\;�b1����첑�![Qv&�-i�V�a�qn�T@�N��g��~��R"e���AY�T�w4�wn�fYpʐ��q8��[��l�wgRqzj{>�KLy�R�lFos�� ���F�
S��=mj����}�������c�E�TP'�Ö:��%O�Fm��컴M\o�j�B�jA��V]�.Y�q1��{ԙ�㘛C9J�5\��^z�MA���\Һ�����"�zm3���f���0/����'�ur1����(�QZ^N�R�	o�ȿ��9Fm�W��ɱB��x,u?b@}T䇓�.5��yV=k�������B���~z�S�z�xoZ��{�q�_,���	_��h?�/�(��d�Q]��N��H��w��@�W�����`Y
qHlm�Χ�����|-'W���/�~+��e'�Bbk�T�di�N�8��`7���qGP��y=��X�*V25Ԍ�z��hv��ڗJV )����y_%�W򻁔{��c��e�*K� `҅m;�f	I.��玐�v�ұ0�	t
5�V�F)N��|x���]g��ccŗX�J
�4a{�|u��_`��n��[C�kVq��E���1M�ͬ����g�۾f�|נ51\#%�E�J� ��=`%x�V䈶�͡%lH9���f��Xm�~Qu#r��uS�"N���	**4�$�U���U�a+xE��i��)<~�d�����>��94\��j.��*W�tLT�b��ļ��y�ZI��i�Y��ZZ㣋�ǎ�9���$�.T;���8�?�ǦyN��;ԩ�"��2sL�~�2C)8���0���O�dl�q����������d.v�Ͱd��Y%��SZf����xq���a��=����5�a��ɋ�Ɲp7l�Ö��m�#�B�&8�a��J�y����9� ��3�>�C�_�T�%E?�w�����C���y�;|���P�oF�70|'`zX�C��0��{e�	�*v<�-!�l�����r�k@�@�b��-\}?	Ů�Dt/�"�>�+}$"B>���*��?����\bf��8��^[�m���,w(����E+u��Z�j�C���j�s'}�l	]4���d)�Q�M��+vo�E��zm�����ټ�RP�ZUc*�o��j�7���������^>����=B�7t.ۤ!�OـA�N��x&��W���{dUTȔG|��2tA��Ω���%'rT����}D�q�G?���f������s���ţ�l{f��$�	�b`V�Ɇſ
�H���OEl|��I��~��%^�4���E��kj!��lW�¯��L�Yw.~P��"Ջћ��x+?F��ڙ������U���@?���ߒԽ�d�lu�l$���x��ԛ\�q�t�pL�MY=˶�h�oH���!��~��?s�ș���3A�.��8GN<)"~�ᐂ���B��;/Xܘ˭%8]1����v��s�fN�k�Lۋ1��,t�d�ul�	9�E�Yz�;�����%���O���8��+\�߳���@^[���o���>uI=�Fǰso���qk�Y����ᐵ��~ֺ��6�G0�hD��i�)߲JW�핲����鏺뮔����N������JW�e
\3�2Ɠoe����o\;�e��^��k~l��c�p|�{�`~!w��x�=n�:��ؓU39��}#Ŗ᦬&�a8#`���M���"�#�%�:�'��FW?̳T�'�2��u�V�B\��B�x%vN���#���˝���c�#Tי��֧�w�j+�1�Po�`Ч."^u����>o���,���^C �����A�߂���'e4��!����Ta�A�o���7Zs�E����>4gt�ߕw�`1��/�L����Ӈw}rCOt �;ݹ�(ڶ­	��g�/~$v��4^�B�/|�yA����̌YC'��*��(c��%WąVJҗ��a2��Ìѫ�y�� �*%�M�Wo�T6M�>�Kҫ�|���k�ȟ���|�|�d�ԧ"�=L���Ӵ��\�Ҧ�*��J����HL��i|����8��Wp�a���6VQ+ߤ��x�Q}�٫=�g�!W�]~6���OHx{��iMķ9�Xjb�� 6Z�	��=N�`f���6�7�Ё#C��x��[���Fas!��eeM�Ճ���"f�����]G#��M�¥u�=�N�%+��[�p���l����x���x��Nή���3���3E�,�tOslwY��i9C�0W�ƕ���n9��)��3|"�5X�f�r�g��&�&p_h�I(_ң�2a����[>"'ߦ3{�-�\��3[b�E�'c݄��/�$�7�ӖN!��ܹ�%��.|k����B�TZ$�n|[Ǩ�s�����+?8�rI���o`���ð@����.��./����j\�V�o�^��F U Z|T�5J��Ҿ8i(nrE�U��Sر�iF*��L3V�@o��nx'ͼ
�I�r�������w\��oS5�ְ�j\7���{\0��{2x�j��������d�cS����Y���˖��� ���r��h��K�X4x���6��H���gv_Z�)=�y)��K�M��ňY=t��0&�kA�U�4.��-�C��ZI��/-r�<'i�H��j3Z���>�sUkQ�9�+���O)�|�.AM�钱�`y��v�ޜ�ce�y�bc?��?7��u�a�*;^X��̪�8<p:̨��z䇵��6���&����x~Ζ�
i`x���lG9�y�&{Uﶮ_mHLS_&���rC��+�9mo]y�-�ih���Z+v�V�%W���V�5e�g�}$��;��h���o��aC�[���q4�����'9>?l����u��)�6���h+��c��A�@G�%b�z�ߴ�o~��Q�"Xi�KC���:DI����G�[Ţ�+Vz0��\����5%#�����J	a�����~I�s��	^nZZ��S��ǻ�Y=>V��O	k6^�V�x{�c/�`F�w:���R�fQ�Q
�'��^�5Z,�{���&�A�r�t9G���ڭ�o���c����~_�m�mb7�І���=�r�ȶ�UK���	���L��ι�/v{9����tl���R���x�)�CO��I3��8*2"ޓϭ�IHB�@�N�a����,�'��ln��%�M��un��m]���.��x�h|��W���\������Z����w���Jr����s���}&2nU'���Xba.7f�'yMo�}�A�*Q&s�tȉ&c�ɍ6)���C���d6�o����]��$K7{�"���{x?3�U��}�����Z�X:�f�s�-�vl����Ih���G�d�;������E$<��QU��F�hv���iީ:0Ġ�}%�V���Q�I��"�5+�x<r���!%n���6��)�S��m(۫z���/A�D��`yyV6�����r,|�ZU'~�q�Q��&��6�ho9�A]�uh�٘���y�G�~��{·'��hT��N�+Nq�,%>,7Uw�hX��׾*�h�����/K�bIS�N3�c�6+p��$'�����7qf�ڐ
�2,�Y�,���3�t�@�飗���߱5�_⸻[��c�'�^2#��O��ܙŜۉ��C�ig��ulr��S�G�r��U������ �/�7G�<n*ͦe�mn���I��^(Xu�r����y�?��j1c��q��3�/?G����<�J�mW��v��q3��R���ё���=�1[�L'��k֦��=�7�\�X@������{���ں����U�BM���O{c�}�e�4!U/)�+J��K7W�8�P�Ҥ�W��#�ZGǪ��o���*��C��&3k�a5ʺ�{)\�9���Yo��PlTY�b��q��;j���mY����<m1w��J�]V�x�i���&-�#q:v�󮿗+����LѢFa����yg»�W�a����b�zpo�
a�����sL空��#�~�l�*n�%%nS��ڧ��5ҬW_*/�_�b��e���Y�L�ъ�X������;�o���ʭ��X��[ԕ�+ej�|���%�/��]7��l�-�g��xQ�����ڙF����ڊi�)>�p?jٺ|�d� �l��v5��)�<vƻ\�g�%q�x}�O��2{V��[��*��N�?'��I׽�F�.�u~3\/�"Լ�M���;�4~�_��܁�G�Ǚ�e]
8U�������5(ܖQ_�n��K��S�� �	��m����"}CЪ���{Cͻ8l'�.W�!�?�*P��r�J�$0�L��ν���`z�g�4+ݑrjԷ�j[�zZ��t�L>���C�o���O��<ـ���NR|&�W�8���%.��<�*�Ok�'q��G���F�@+�t�3�80�������Һ���^��#ލ%��5�M�#�f�#ّ)9`�"^�&�b/%�_ǻcb�6�I���d�w`iRK♨"7*B[���D��Ԇ�����nS�7�~�ws�j-����i}ye�%oP:�Cx�rpu_������W�q��`�ֺ�wf>O8�ݫo@²MT�%9Y�H����������O��\�4S���?_�:p�����#N3����-"#��i,5շ5����rJi�����+T�~۠t�P]�F�m��#�i����H�v/�$wk	���5R�aў�t[�J�tnY%\�ZM�xPO�+"�GV��#1�O�{*�t���V�w8"�6�N~�½*���L��n��~Qʇ�=��/��+����E�lED7MA@E����HiҔ� t!���H�"�R���t����IK-@��I����������̚Y�y��Ye�;�k5_˞�lU����f�xw��K�S��Ss�R#�Pr�'��?�yfD_B��Ӥ���W�h��6l�1̹>U�V9�v{���q��d��s�X$[p&[�w�^��I'��Kt.Ű������T�����_m��!á�5q��?.���w��1u@���ɻ��ppiie��T�qԖ��p��
 ��B/J~TvW���������7v�b���>�<�!{G>N�$�z�L��"Q���m��z^h:�+�Z_�ĕ����L����s��w�X�lŞŵ�oRU68�}M��'l��p;5e����HZC�ꡨ�wo�II���߾��`�����l�i�+���Ԡ#'(�e�*H0S��BJ�U�^�B�}�*��5�i�,�VQ�B��	9t�|�a;����S)��DK��+5�h�~�X��*�~��RJn���U.oZ�Q�puf'�M�b�ێ+[`߉?pM1	]E6����c�"{����_���+��r��u.� �I��^���RI��öe�<�>`�M���L��WI��է���#0������Ƹ��hڴ��޻Fݮo��M�ě��FZ���0='��M�:&D�&܀=<5_ڼ���F@zZM���]�QG�
S�q;4}W�`J�h[*��Y�g�U5�ߊX���o�9�xX��v9QpA~��x�	����:�	�FQVtu��[�73&^5�Z�l�����6Ӎ��6���/|\�@I�'�����.��9==���hD��9}rXQ�p4|�<�GP;��ꥎ�ʹ��')fW�{��ejNl��+s#e��fi?�&/��׸(
쾊Vs����g�Lǭg�xOՒ�Ƨ�-�_�y:C���@rn�IMy	��b���_��l��3T�>\4bl}wl��6��K�@,����"�0aO��&GV��`�z_��o��⼯��G{���V�6��m�v�s( �Æ���d�k�Orzw�;M��.h(���x�ד/d��]]�$����ċ#Y�1]�¾�tuo�mG�Р$Q��i�n�u�R��&ϡ^�LJ��ަP��m�SG'�~��p߽�j_}tX#�׎�e�kq�/�>^�#����?ȉڛ������Y���:^��|^Ò8����[���0�vsa��=��˭�5����W����D^��Vu!]�u������V��V�|-&.�a�+>�d���0�S	#�_V��ǭ�=<E;�8��{�ڄ}*�����@���}-��̮qS�D�Hb𜪜��;��x�<�u�1��ݜژi���ƈ@A8����fSy~�v�p�m������͟�8V��K���'08�hDl�(~ *c/LR�m-�x/���?%Yi�/�+�[����3ea�Fz���'yAI�%�Uy�qd�^	N0��IU�4h�>dz��(x����.�7�R��L��L� ��Z}7g������=m4��wZ�S��)-|�����+4%+?QMNv�ݺ�~ks�2�PD
y��	i١x��ZV�!s;�>�����ow%���#֫k�F�J��&k�Je�<ax[9h����e�̏�U�h -A8,��H3�M�'�����9U�<<ʵ������ց��q4��#�zN��io�r�@}ї��͈:kep�a-�n#xo�U�\���;��&י�J�,���9���N
NHPe$l]�o�7#�sy�ͪ`~�ڬ[��c�"o-}!��p���+�/�wKT����/��)�oNT�y��>qR���c;z��LWܱ�	���.�`%{�+�F�̼7�!k��eGa\wa��u�x��"�/���f��_��5\f�wJ��������	���擯�{(ι��u�o	�`;x��v��Q��&�?"�7�p�� ����;�,�a����o�aU��~ū�p��v\9,�pr{�P e��������������@�
��O����i��E�{o{�����޶Y<���\��G���W=����F��Ɔ���좃���A}�°U���́~����������sϊ~'������$$�@Y�L�:=��K'���hI>��֎2��ܶ/)k�\�td�����P/��}H?������d�`��q<7���i1�=r&/x��m[N<�.v隩Ʋ�\?��\E؍}�Ƹ��VX.
����&�F+g�cX<��0�.��g'r-C�;�X��yH۞v2�;��{�S,8t�p���iwW�5�]Of%`�<�J'պ�D�n`A�>\�SVBe�Ezv�xzC�:	y��˿���I��D��!����p�S �+��N��:��L�
�RbK�}�h#��:[8R�S-$��f?y�� Jlsykȋ��^��[��2l<�N��K{�=T��h��y�4eyV]+��1�^w�D[r Vz��W���ԽO�l������Q�	�[���4�� .,�뵺[.��r`D��@z�����w5����G����[v��ȩ��=�^Gv(����h��
��x�[�B��'��>��?���7/��'���ķxq#�^��)$���Ǉ��eM��F���t�OE%z-��iik� �K������|�Pj�C�۞�tTi����|��K!�2�V��\}��2X�
��.��f���l�5����/"�S����Ŗ��䫍C�OL�&�S���n�@%��hprʞCi5�
�����_l�����`�X�D1��c���e��a�s٦�~����+CYv�)�[�����ȹ@0I�]$u��B�Q.�e�g!�Gfݡ,*>sJS��[MR�?	P�Z�i@�(��+ �+�:k g�.|A�p��h���L��wyM^����e�P(��C��߿����5����],�Ŵ���0�ܢ�-���9�˟���X� ���Si��J|<�:+]��X��[��FU�=���ر���aS��6 �������8c@��S�Im~t��u>bXh8��iJ�px��y}����T��v�,Dę�1x�l�o{���r49���V�h5�q���W�G�d���h�1���9m�j�g��g˒����7$m*����n}эZ��z'�3�Hݞ�j�	%��M�ZW[�F.�^��]�"���b�yAU�V�w�nQ_���1�~�!�q����W����8��j�s���J�f]u=� Lϗ���Ӟ�za�j��k�m���MZ�N�y�zc�]"H[�=�gg�`�t?�mR_^g	��)�������ŇX�D}���TV}�K�NèO�u�ަQ�l��:�T���R�4)��~f��s�qߝ�L��T7{:���P{��Q_��mi����H���%?*HBb.9"}_{[z�>��S���-3n��%'������F�I�5�BJa���?�7)�����8�������+��e��)���{��5frk��]è����i+�R�w���ߡ���7��G�\']}��*��� ����sI��S��\H��(�h���xF���XSW�rnb�n����*r��FBE11t-�q#N���T�S�0ջ�s���I�֟��X��G������Xy�����['�?�s������QH�?��jae���d�
��I����ZT~Lߣ��:P_Em*��-q���[�0�~������V%L���,Lb��e��5`@��Z�  _,V����es]@h$%Z8Z������n>���u߲@-=�L~:r�>��^�w~�j.Ǫ����P�xݩ��z��r[9`����=Y�/Ԅ������s��R��;l�>��7n�2&ٖMJ�����v����?N<�}��SM�/@B���X�q
�]���m���?�㷰�A?M\Q�_e*ab��; ���޽?C��{�)�:낲�$G>�W�V�]���+]�����hkÌT�M��,��M�����z���dC� #Q�IE���\��K<���U1�S���v���>�<����r2���D'v�
{cO;=Ջ�ihD
 �m�p��"g � 
m�ý����bT��7X�뜭=�a����F.&7<�;E����� (�y;�v���^�嵫�[fM�]Wc1v�| q��د�ɹ���\����ɾ��>���Z�%�+��ޏ�i�{\j�zW���+}Uj����+yӞsk���8���D�g�m�7��vz�����
�Ș����'zn��ՁV�^t�c(<F+-l�6:z�LE}�`T�t��0���#� ~q�����dv���w�s4�iF6�R������1�������/q))EVN� ��ml):�Q�B3-!ة.��ytC�Z�rg�����n6@:/qt>3�<��2'bN�2YG]6A��I��Ӕ�=T_����[�
�S�m�v�W	�ׄo�3��ز���n�o��̼�z��a�%�{x�X �3YSw�RX���Rw2�jp��y_c��/~y$/$���b���D��\���O���v=��5���ȕb���G��:�}��[3v�5Ee���)8_�ANT��c����x]}��Q��r1G���b��q2a5�nJH��Ij>K�d�m���<��ރ!ݘ�ї=V�¹��^��DU���1��P^'�:5	��0_Y<#�\z��b�E�ؖ2�T"}Y %>��9�A{ #@N�]��r�) ��Z0�n�,��ut�G�]10���v/���wj�W?;C/V�]pEK!iQ�ƀ��{{y<�! J�0���ץR���=�eY��>��U+k'"-~폊�����Q��F���X)yٳ���)����vM]��C�Ťl�+F��K�a����N�|E_A����kˣ��Qo��Ů��[��X �L]�45IO����A_r�R�`�d���,1�����}���e׬Qצ΃<?���B�s��_S-�KS�kQ��sQ/U�� ���osե��T&"p��\ْ����0����/�ڋh�Ɨ�[�;Ƌ�MK*e�B���� ��X(�\;ޠZ�����V:Dt�6�ЗB�`w�Ǹ�ܸ���b�ݪ��ҢW>d��\:#_T�^�$���CW77߾�K5�stU�qX3Jt-e F����\]������Q���5;^��f5n�s;ݺ�<����q=��p��z%4ڗ�E8:�̇�y���6�<9�i��o�=��=t>��)dw{�fb�~]Q����i�'L���9Β.^��6tҀ���i?�ۢ\�ꥮ��b��:S?���u�����e�"�?��QH�i�V�&?r����@�����[�t�EϪ�C���{+upr�m��j�$qԲ+�\��T��ѫUaV����Z��F���m�%85�j�Ar��N�,������lbWϐ	�\�o�\e������dV6ՠ�ѽkӔ�]^��Ւ���}�x���K����}6P�CwNP���gv7�d;q�Nz����3�^�����^���=/Ʒz�"��Q�]��t�a�Qu_2�/W��� ��S8�t�Z�����MT%z�:/����4�:�/J&�Tb����TLjbq�^o(����⥕�u���<lF?���8Ƭ�́�1gUMR�/�T�h�Ű���������d��T�P�����k����\��5ٺ:�[�DC���R���Ґ~����YݱGS����跴�x1q�N�-�e�00a�jh�;�6L�3��iO� ��/���eO�E���U^c����L�[H�պ+ͩ5������3O������ئ���x��u�G^�@����$��"�g���+!Eg��g~�{��%2���>q���L��6��RN���臼҂FOb���Ҽ>�P� 6�oE2ʘ�OST>y�~�Y_"��g瓕+o� �������w~�R���{\295��~��{d��"j��b�l̂`�����{:n���b�BJ�;��<�+�������0����=@F>:&dce��y:�=�� �����#��l�e��8s��4����n\�!0����1�OP���Ě�Z�I�� @�;,U�`_Ҥ�i%��4�n+?�����um1o�/��A>c�Jݩ�<1h][����wL�l�A�����i�[@���pj���e��:ݨ����逄�K*��ѥ�-�ŹۣK�c�L��,dePjz��:�<}�qA��3dk%�k��U�|��'���������,N��o����\T��j^���;�E<2�n1+�I�P!	�t��6%��5O3�C�SY��n.���L�m`�������g��5�?1I����{�J��OG�l�LH&���2i�$����#~Û|��N�ig~$��[k�u�A� �)d�e Q��0l8��CbI}μ�˞m-'O�^�u3����W	��:#C��y7x���fW� ��{�U�Qޫ;R:Փ�C�H�Α��4D��T��y84wNܞy�>nXY��q��}Ss:)@��})�A��S�*�P�.o\g�ίH w���t�����)������c m �b#��QMFE
��SD�p���D[/�.��
��;m*���şl��lWM�[����̓J��E�S���@\�נ������b�O�uEV�0�q����A�g�u�.J<g��v��Q����r3 1m(S���?&CO?\Q���9�XQL�×�A�FL µ�P��D���A ��t�6y>�������!>Z�%tl�uZ"��ȡ�ݖ췊��8Rw�_�n�Q�F-$3/j��Q�|�i�3c8nL�|�o�.�;�Yo�f�g�UY�� ��� �?q�9���P��E �,T��t��)��{�Q�ŪX ����v4�)�@����%�H
/�%o<�N"ҧ��L�_�w�!���^�V�چzca��E�E��e�;��N:��}΀����ID�ZW�t�s=ڒ՟B����At���{~�� X���;�Tϧ��r��|�P�5e�WY��В�(UJ�so$�+�?H�ۍwHeu����?���3�bũ����w��XpNl����4��/ʇn�#�B�r#�,��c���y4z�'i��De��ڐ+I>��@��8���7t���#��y����n�����y-��/q��?ӧkۉi!��'��,����|����'z��1w?�bˏ�!�@7f|(JW�m\��3I'w�)Y	="����{6�S��u_0�	�l2l �V�J~��M�%��D����N]�c>z�0�������#��x/R���|��;ë;wXy���;>�]��/5��;�Z@!�������qw�?1�۞1m�Gv c:�B\1%���A7��;i����u
c.�J��=�6�4#��3��|���=Y'0���E�n��y��Rm�*�s�U��:?�dlc&��սIk	��G�g�k25z#�}Or�1o$�D�uj�`�zݳ9�#Pz5�O�+A�?�r����'�-om����ܭ�R_�T@��nRAj��ቃl_�N���*�H��:�*���h$I5���Z܄j�ݾa;L���~׌�|/m\=~��ř���$�w��?;��|�3))f=,���|� ��$�R���	��Ŧ�<)��Z#���&H��2��2O��ϖ:aYZ /ۣ��.���8���%Fݾ�	�=nD�P��'�}�F�.#?�
���<�_=w`��b5㌟�`|��Zjd���S��y ȒV��B>���-/�e��|8���V)Ms�	�8���{}
�� �b���ɉD]���ĕ$�y�*��b$��q�-�:�����Se�RV,E�Z�/�xr���	�*��EL8u�^|�q��k@����X�z��N"���|�vWϱ ��h��JN�m���|L��\���M�d���3:�N��8�МO��J/��	�a��K�t�7�;ޠ��]V��]�@$0:��t�\-�3q��҄��l�K���V��u}q}��ifk l�'c��� �67��W.��*��
 ��#^���@~&����_�l�.9_=W�Ϗ]��(v�MƟFw���7x��Ӆ�:��MNֹDO�3ҧ�_���J	���������$�F:�#�q����wY0��TwaA��[ͦ�w ����Ѵ=�C�ĀףS�DȌ�������"����!I�]�,�s&��L�VT�qJ�-*?��Cz�t �mN��m�O�v���^�:&�zk�8c�a �	g-y���d��P0*]� ��t� ��$���8�����	�����S���!W4	���>��&���m�nL�_����w��*_Ͻ���r�����O	^� ���U�$�f1 �ĝ��Mب���T�{�?:0�aFω���l��B7hF
MF��foS��k�_<�X0��i��N�0�fv:q	P>L�&��{};���d �'�=��6��]�SZ�T�v�DɺgܦA� �`n�������=3���iҧ�8����M�V�{U��?�?��N�dR��j���x��N��Hu��c+ ��N{� ��ͤ����Jfrm���xm��Υ�J_5��+q6�`�ܾԊs��4>�����G��`dn���%�l:'�#��RO���BK���%:π�/7��&Yf�%2�1_�b�<n~�X}���0M7�\<��4+�D������Ĭ���T�ȕ�$i�7NAݣ��u��ؑ�����bzap�&��@����<�M.����W΄p��JyY�tJ�jA1^����諞�|����:8xJA@�PKC��{��Y�5�:�V�)H&L�c��R�F��h��2��f�bm�&�
�IEcK�ޜ��Q�f�QqˤIη@`xm�V:�ۗ���Ur5�=��]�B�W�D�;P٤G+��0LR\�����Ӿ��U�F�"���q�� a��r���ssD8���jY�T��Ԫh%�Gq`�ol�K��{�� Z�ۨW��0e��»jH"y����	�V�K�}O#O��s�Q�$.��[
I��`�t���`��x�&�U�븱��
YK�"��佟P�Ƈ��è2�:��������\uZ
%��5.f�_��%Ӿ޿\4��9�ښ�Rp���(�3�`�Cx�R�;�/������85Xh�n�ׯ�~!WhdIjM��@�I���L��o��{c5�����b�x���t茯�V|�j�~�{�]O��L�35�
��S��@����v=^�HKG��E�PS�']�7���\�����_U�vfb���r�Щ�ރ^���i��"jυ�AyS�qe���|6��E�p_�i
������6�N�X	Y�� @��q��h0l?�W�}���w�IT@�&d��SX^+�&�z��~������5���J���sߡ�����iT���Ҳ��h�[g��sJ�[��Y����?:ճ7�|4y����>�ܡ/T�����!n�Q�3� P*t�D^�NA�6�51@���Z�(񥈖��DIp;N^���H�j1�Qq�ᰙȽ&���-�������=D�4�,���hء2�����k��q�y8�xb�X�տ:��*??�k2v�� �C����ӻ�;V1�SDjng��Z���qy�#l����4��O� �j4*a��4��}zuMf�@.��j��5#����5(,�4w6'�A�����P;������	���|O��Qت�J�'����{���Mu�S��;s���1���o|��ou�瞥�S X��PH^��Lڄ�q�������}�V��_8���2@��r#��·����9�(�q&�m W��iq������}�����%v1*Q��M
��b�/�V#�_�ۗh�)%|�J��k\���q=*�X���)�iO߀��������/����Kҗ�G�����뗨U��x�&���i�c�|�$|=Bܷ��2����ntN��C�+�����v��6B&���k�A؝&ai���Ϸ��Bs{o�=��M�/%��T2*�\��L�,�f��xZm�]J����-)����� բ����k< �t�/Jfmפ������>o!r������j��:\)gv`z��ִ���毳m�w]�t�N�8�a�c�A�k�����ܥ3.� �`Ϯ��C���%qL�T4���)�pPy+#�����J�{������~��{�E���u�&�<,��_�����~���k&�Kƶ�q�U�=�Ә�����h�n���O-��y�pl���m�`j��d0�����l۷��̨���pkfR�������[o���vj S��W�PW��[�o�q�(�͵
x�����!��|�7�z�x��d����/��M���RDn�'Q�{��-'k����餚����K�f<W�����(L|j��VuoI/�W��)#�sj;Œ}CaN�b��|�������@uZ��t�n+V��vj���jy�!2��㸫�3C��++��\�A��v9�"28�f4r�%�����d�����y��Dr�R�n-�r�a�Y=��-��G�����{�����-�����Ƒ�n�)��vn%�{�y���pcQ���8�mp6#��[܋,a%�|}�Q�
:8�з5�����h����4�(YC>�����x9C��I~�V���&@(Z<zi��&�w<z+&A���b��EG��Ԁ���	mY�p�|�����d�格�$۽Ch+��p.U�xs��U�r�!�:��k�NY��f�Y^�4�]�/����|�솪��;g��8X����mY|`���w:�]L�屣�typ����f��-�T���}�	�|][�v�A�}a���pWy���q���,;�������c����f�9u��������9�yı5�5ֺ׽%�?-\�4�u(�~о�[�]����^F��>�����+�1U����~��PuW{�����݋>��S<-^���l,�	�:��C*�=�`beۤ���K��>Dԋ���Ϛ	2�<���ߔ��7���?�)QVY�)�P�ز'���^���/�#�
A��7{��J��1m���06Ԧ��d�e˨���&���gV�\�YoapZ�8�]d���C�.�� G��=?�7��;ݓo�x�>�^2O�\��� X�3w�~����t�d�n��A���I�M�!;�K��C�*onnl2��U�sի�?��S(
p	� <�̮r>��ً��L�ں�X?�c�a���7��uT|׏�!s�Ж��u[�9ŵB
������H�꾑햾~E�����j�ثv)�Ӵ�=Y'X�)�+,-&�ӏ�Пj%w����ױ��֮��_�`l��:Υ�<y�5l�z��k
���z%��P���<$)�m�ײ�s[i߮d�^?���27���hz��Q����Z�7H�A���
��[v�b��F�满e��9%V0M#㭒����UK�g4/���0#���a��Oo�*�w��9��*������{,W6�X��0{�&=I�0����MK�{<���ז���s�/F�w�zva�3J���u>&u%#�f'��%w6	<�}���%���e�~�⺂���%�
��O�SP���oAP��RǍ��]��*Jݭ,[>�o�d�P���yW�F�*ڌ��
y-�`�pc����z��zj��V/0X��Xݤ�$>�q.'D�a�-��Q�'���ѣ�N��}�Q����X�l�6C�����r�1_�ɢʒJ� 5/�1#�R[gL�G��G}?s�ʝT�I��ۨJ{L�l͂-4T�~�glee��Y��bp9YYJ��K��A��@�i0�^�q�UZW�#�W�.�jP*�dd����������5K*���
�D�E�����i���75��+Q�ښ�G�\��OўA&�{CU0g�+xk?���Pn�g|宲�pA1'���=�)���#Fw��;4y!Yzf�����J8{���IMjh�������ǭgP6�CmY7�(��H:v�-�:��e�9�
�f��,p�2�!�D�:����f�ú�q�1a���B/���KAq�\��/jL;����K󰆻	��З�.�'����ߦ�rT��9�M�r�N6g����ʑr����U��ʲF��p��Dq~�6�3�,Rpg �S	o��#�PSL�3���%%��r��+�I��!�}
$�p:A�Ŀ��e���[[�+²LM��� ��u"i7��^��v5���q�2�r��G>�w�ԑ��Nє��2���\�ocr���u���M��}�k�+	��-Չ�]&�Q/\��pVaH���[h�s2#/W�"ȃ�gj2�<����g9.��i�w�9����g('�\o˛�p�}��δAe�0m�f"Vqq�g�Ⱦ�Ϲ��btm�Yb�p2��a��������y&IuL����X����tjx��Us (�ck�~#%>�VX���4A��y���C�c���o>!d((�:$���O=e���n[D���^�Uu~p
d�m�����~�B�ԕ:��Ć_�����D�����B)=��Z�sj���7���ԫ
�$��rX9��Ww! �{z2��Y�h�nI���.�R�����@J����=�ڣ���_v�QIu��ab��
 �C�K�F��5�QG7�Ӻ�F��0���L�M�;�����{����NcM�L���Wy>$Vjs�R�2$�yFь�z�3ۢ �g*�w  9��k�)�G�n�tx��ٷ4�)�K�K����:�2�J67��$"���孫c��dA_�@����D��\O�����ΣF�J���k���O�m~@L�>�%�K aRnH�[�V��m[����RŐ�>si��.�(@#�;'�x ≣�o�Uq�[��L4�_�TF�r�G�½u���Q��9�R���U"TBnw`d��ڎ6Qd�5�����gI�¼>�,��g�]]����	������" �HYE��z� ޶z�{ǁMXL��ငy��ðՋ�z1��;�)��Q���Z��޴���EY���r��8D�'#7�Ł{���&��AZ��gv�F���r�?�*\�N�7X[is�j��V±NΔ�5Y���vP()�%1�yn�� oH#���z���feԳ���Y�^� ��� ۮ~[&M>��v�2Zmaa�Z@(�L��_3����' �աA!9.^Q���B��������abط��MJ=?ڬ�O ���������D�s7������� r~�2N��
q���t�����^^��'�G>Gw0_�,{�W,\Sd��c���r#%�����Cv*�F�����1��v�����P;�C�{�_ħ�ӿ��"0�>�C��,@ya��h���	����V����C�Y��E�_
��:�WZ��O[��}��j'A��!o�l{%{*<m������q����*`̗:�&6��F9x��Bq�QnwsDj�KddwrA}{	z�l�31���de?zo� �1��_�9(���u�*�铞��N�� ���ji/�1ҽ��^�����Q�by�Ai57m)��RA�#���@�$&]���iM}v��Җb�U>i��=���tٟ��_����%���1SF��VO-Ŏ�5Q������5��9t�Dk�)�����9�ٳ.i?@�GJ��xY����N��W���@2�j]��ۮ�(ߧ�`��1a�ӿ�}�����Ж�P��M�6��2Q�<ۮ�
oG÷5�$������W�Do�#��܋z�����f�%id�����n��R�D���ͣٲ�`�e���V�G�^�GH��B�M����BIkS*�3�/��^z��~��b<9X�a�j��ܨEo=��|T���D�Z�X�-��WA-�7�g#�W�AG�p_@6U&��]���)���c�����3:�W�gj�ꏱ���8n.��@�㣍7L�_�k�6�[�"*��Lo �t��ӻ\1/W~H	���U ��/�I��Y�.�P�M��Hy<˼��'n�Q�y�İē�;��#�ӄ�qq`WV����S�j�ni�����6����lW�djyD�����":_���_P�"P����W���"�n_U�oG������Y���J?ԧ���WM�?Z��F����n���X����ϴnƌ�Z���w�:�_���|BfnaXsR�h,�th����
��I�n  'e�,<u��;N�/6��Rp��@����w��}��z���)�K��oj��;���#�a��?�%���$�klh��G��Tvފ|�Q�sA<��9���à۟��VKKU�b�z�4{,�C�JR� ���v'x��2����8��UnƬ(Ȉ|�V�_��nM���'�;-��D/�}�:7��ƨ�Ĭ%�H����G�&��6/'�m����М�?9�3��;�ێ:3�!�+
������so��0�EћnvN��Ȧ���� {��_ߪF�K��+|@*��(�/�#�7Zv-�^�w���X/��ĘQ}D���|磂�g�?���r�e.R�*�]b�#�1����uZc<�-cX3!��k�N���:�E�-(�˼9��O�K5�c�O!�
�(��+��K�/		!����^K%H$k�L38�_[gyx�f�exO#i�u��� \��5�A��|�N;�fY�ؓI�i'�GL��9�+Č�bӼ9����(��7�a	�04ꀘ���"�B�����&|�`7����k!#�������I~����1T6�0� 8��/� a��!畊r����&�m];�#�O��

�o��#��U�S���k�	K�^��E^%?i��]gA�pu��;$GjQ�/"�3�����y�v�
���?��M\��-�{=
y�l$É���Q�=�H�z�`%��v
(E�w���"R3�
�������:�M�N/�p�q��N['���S�f�&HK� �Q��낍�C����*l�{�cc�Pu3�}~}�V�bʴA�25��+Y�y�\k�����T%������j><�������3�	7�����#�k�곎>ĥ���D��;=�v��і��D&|��@��3
w��g�]���K�7+m7���NWg�4f'Р������ƺ�Lr/�td��|�/q�����=�\�	u���?�J�����k��虑���������M��ݝ�HY��57@�����.������I�z�����͊2���N��I��2s����*�̯&��B{����AAh9�U6#Iw�>NԻ�� ��+�OZt�A����;���t��u$_����u�tu#W�(�:g�&&&����֠��(�����������iz��W�b�����P�� �w�Xg�)<U�hr���H��J"���q�)����uu��۟[�+��0�K�z��̦z}��ȡM��+T�Սl(�~-Թ�i����<� 8(&���RW4����0���"����*��S���y��;��;�&3v-o+
�� L�@�;�)�a�@(�$lY������SY�c�~6���.�~���~���2	�=����+0��l�d�4��P_^�-���HQ�7��(U��&��f49vu�LK��W��cM>`�w
��իA�_T�6����YI�X�-Q��_ãװ� ��?
3M���r�^'�(g�{MW{[TPW�kj:\*okV\/]�p�
�!���ffl��^/��K)E�
xRo�,�o0a��(m�g�o�y���C,�W���++#�4���Dۛ�K�@��nb�Ǔ���	�"GhW+��)��N�hjjv%���Vi��Iۯݦ�f��H�[)�q�Ë�;J�p�����q,@�v�=����r�-F�͵kH��6I6�iI�������wi��w$��Ju��uW|�p;l��2�l�,[5kF�1�;�t�	�j�{:՘�[���6�%��}��)c%g�2t���b SU�ԉXW;�_j[��a͜�/��������qż��F�t'�{N��k$K��v'K��z/&��z:F8�2
�gSԋU�l�X%��:
��9=>�.�����Z�v�ƪ��#L����w�[�J\��Ϊh$���4f���)��@�%�ޣB�Pe�11g�w��W���֝H|W��\A:d�c2_�������}Ǻ7�%SGEE�����p��/�i�"�/$��hA�k���h��?䟯�����J����3k����4���y���G�q�%�V�q����M�O�B�$R0\xnY~|��V�/"is��CDm�o�-Z�6e��]�F¥]�,Gk8OH��x�?MI�Ϧ�+w���V!X�}�F�VrrQC:Za���7M��,��9����Mq�I�p*����Q�f�����C�k����v�ׯ\%��ZTtڡ��o�Ł���4V��P���x\=�9#����޸���*����Q���|�7�8��	<O��R���q6bhty೰�bW�\NNN�������!;����r��ol�����i���|�wp������P ���6=�R˙ѧ������=�M�@�|$ϐ$kO���o���D�_�s8��}T�VO(���ymm�&�Q�,�1t�%&)����q������+����q�ʡ�í^N�;�}k�c]�z��Kl�/?�ѡ�3�0<��p�NGGw8��c[-vV�O��F󩧀�j�6�Wp���p Q�S�j�|����&��
a���qq8}P��U�Q����Q\^jo�/r���r�
:�7�G�k��#�4)lg��K���������D(�����0Z`���{):2}{E0�Q	�
9V-�^�v�\���@up���)� ������iv,���+R>9�*:8�?ޯDW��cQ-�}ӂS,����il����9Y%�k����� ��i�,��$4 �������e;�R�y�#8=��R]II�?aAٖ~��&I��$⟯7�[7�����o��~q<�]�����'��Ä���n�T���������Fy�zCC��\{Ϩx �eklϟ�9 }ߪ8/�47Эu%�ċ���,]��YI�AUYQcCmr�3�i���ђ����8�)���]�RW�2��W�����l�7� \��b��%
���% w!G	�ֈ��/ӽuf�Z	52w��E��y݀��X��"{I3Vx;U���O����O��B"�ظfdH�ظ�a���d�%X��O��>�G5]�LA9�;$#^�@��h��OOc�ӽ��a�>���|�]f?�@m ��;,�O_�z�{�ϰ)
2o��ڤ�Ǚ���/,�].��rj���}�""t�FP�W��׎^	��޽��4��xBe�[��9C��Z��������R���z��sb��/��LKTU����yN{��.��k&I���Q���:���^��tO@MO��������3�7)qw��Q���c��q�[W��QA0��P���@�II���AA@I�\�X�AJ�kw�]jYX��"��ǟ:;��s�����{f�v.�Ͳo`��	o �����t��?ذk6`Lp�s�a�	�q}�=zQs�`A�K�P�%�pg}M�_x��������1;�孡�"Յ�&''K'>Q%��>�q_�5�O��}E�ʅz���2l�D�ҟ9��@�Ϋ�R�� Whs$���K�p��5浸�5��~�~���)��R/�?��Zoe#�\�x�����P Y����_��_,֐��Tu�<�<1����b�b5��w�M{� e���y�����>?m)cDu��������@+�%l����'��~�G���8U9���D�Ŏo�ష�d4�C~U]��BRR�8j��y�V��H���Ѹ��j=y�.yPa��WD�+ �Vyp��_�x-5k߮��1��'gc���?�w+���ϯZ^��`gD��$@d�0��S.\����g\\\�D�r[�A�vvvl�Q�M�<���߾���'$)���<�e[6�C�%�}�e�۟xM�pS�{ȵ���3��*�4�4��|>K�w�� &R����?�_@&�	0ɉ�+��y��f~��OkkK^�] �'�9���y�;�:#����@�уW��m�ʟ�ߣ�P����,yf))��S���`sR���=Q9:o�bj�w�i�.���12�hW�v�/  �Ρ[�C.���H;���>y3�?&&��"��%�\FW�sõ���HSΓ�z?%�~���zѽ����)	Q�B�3��K���|ɪ���iڵ�5�{r ��,���!J�B�&|n�O��������meŲ솽��GXf�{EU���zDb�H��V��7�0K�a�jtU��m��h��4R،y����uqII�j�zd)A�_د�ܿ-���!��:��U���ɩ����������q&���է�6�$�J�_�.��k5i�6��c��GT@�e�=��!���_t��n@t\f"m0F�V��+c����ش��)**�����W��;k +������gq�~
K5n�L��O�x�P�)4dԪFXdA^�fW�.C#J��s�{�Y��GwU�?�u�5@=%�&r��ִ�~��y�����ަ���i Q�������<��MO×�`
.N-ē��Z���	�Z֧m���+B=а��+%��cƮS*wZ췱8��gpX[๏)].l�ۑ�EF��P1C.d)�F�]�g&y��Y��[��-+���ɭ�;���a[��9����N�֦4J�p4��g[��y�h.}�P�ŖT���r���m�������m,�_P�����U�{S��#1�D�o�he#|��c��d-ϩ���c��Ϗjll|������c�cp�z�c��L��w�[�5(������ڜU�鱖�n�2Ɨ��l���À��� �x͓eUU	@������f�76k���/�b=��S�K%O��l��v�gP�&���_Q�������4��$֦�Ԃ��Dv�sAec��
�$��(��5Ԇ.FvXhX�i���V�n-�c3�y��v���ਠ"���^3@j��l��rQg(�p�_b�[�On-�U��l�"44�qCH��m7�b�Ԧ��;�����8���cx�3-k���P�6.���7�|��4�����\uϹp��1d.�G�l5{�2Ƣ�7��=�P4ⱬYk����!��J��(�d��XP�s?C�vlRJZ:%+��l�tk���M�����y"���Zʳs�$e��#&k���($ �Ht��yQah�0���vxDC �1좕 I��+�p�y�ѻ�T]���({�߻�ml��F����sm�rr�ʲ��~,tk>%�>Fq6�g�z�&y��Ӫ��Eo�<rc���%BmƖ�����+J=�w��j2�Dw[C����÷��J7{���7�v6�U����?ۋ�5�el�б��P�Z����� :��}S������JD?�$��a:2�GB��ϱ:�|��LnQ�(�?�۶�Рur1'?;e��`�v"�W�؂�KG���i���4_&���	4��s{pO�"��ō96&� �*�ީ���bl7J#��c^5�u�8��HS�d�dj��8��S�,y������H�ӓ&��2����>�[���?�R[D�0?f�)#�F�І��ޜh�&�5��-ʑ��ꟲ=�=�uݐU����`�5�M�8��+P6?�F5`����ݽ2ii�)l�c�ptz��h�+ύ�o"�q��y@#�C��<�l6���_��m_�����JE������_��G�Te��<�()Ȝ�|W������J%ZZ�&����y�\�|��%�^Y^Ԏ]9�]������j��u�B��WP�6�ߍ�v�j ��q5O��J߶�z���'����~ ��_r�+ʞК��au�'�7��n=f��Q�Q~5�4�����!H�J �ť@��Ξߙ�9��=x��E��aN:���G/�_|�?���r������ƚ��ӯ��x�? �5�6@�)���������E ���_U�z�`BLH5��N(\���=�1�[$�����^�
���O��'	Znϭ���H�s:�? f�z^r}:@��|�ia���vns< �sb�h�}��M��ߣ�m�P �^
�ʧ�9��=y�~��ǧ6��h���X��S��T�F|��|1�W߅�z�F@��7�$����t��[�ʽ�֣26Wh�;Z�=����,?��_���*c}���t��8�����"�mY(��%N��X�ɉٺ��>$$DAE%
v�o7?�<,�y���LST��߫�u��?��"��a::���C
�O��rx`6s�45o���v��rG�|��ծ�n��'`EѲ�pѳ%C�s<ǟ~2�2�-�-�9agz�:'[�us�J��I:���<5ގK�n�!tP	"~��U�g�訞�ccc�⣏Q���!�q�Y7['U7Jp��(tn��S���,�r�>�,Ot�Xy��-����Z�;.[��M'1�=G�비�Ը�~1������g�k���ﺌ��h]k���mM�!��AAU���ӵV���#w(�Ӓ5[V�yM#Z���!�-t�J�|s��[j~�屋���'	Y��%B�R���{���oU?Ӹ��R�\8�ö�E �I�o�ɿ�:Jz�%2>nd��������b �����G�l�o?*;�g�3���
��g�;��<�s��O��.���2�8���0Z��0O��]u|+�_֒�s&�:��.�+1�?��ɪ?j� ���T��=����Q�kӉ�m�h�k�X>��ϬAd���*��G��Gq��n5k9@��O�Ω�ֲsR3���Sg���&�!'O�}�{p��+����o
k��L�&@o�8;J;\���9sxy8U�
7k������iXTS�@x�%I[���O�����]˕V*��$�����ʙ���h�*%���c?>aN �0�qq*�9�oǟ��0Nv-v�,����k�����_c���^�L��YUS���M{�n[GOӭ

���h��_�����ߩ��lؗ�%z�=���z���U��Im�j�&�ZkA��AR�e��R�E�9<�z��P�HH��Z�w�4�5T/�����s��bA�#7�~��uyg��e�|�c����%,�tTp�����f����ݴ�. �_�㸨�z�uYڌt�O%�Yc��F�����T�`d?��nS�|"i�*�8���3̡��a4�`����/�}B�j��weky���b{��g�4��������i���FY��b� ��x�үY�o�����M>�"���^��ӾX�������0�/SHg��棴2d�rm~!	�S�0��bЮ����¾�;��N�s�E�ϟ|5;Y����r��ng[�y��m58����'g����%�J��@-�e����{{����;jX�ش(����D��s>��C�A��wiܲ�	�N��sd'?�v����q��Q������aO,�� x����-�Avn�D�J�-T¡=6t��Ö��-ulD�t�<b\P�z����w�(V��~�����|�٠F���َ
�&Z�a�k���o��/4�YO����(�0#�ҕX�z�.OAV�D�>�T��\��i�λ7�o3������#���L_�=j�ۆ��.�����c��U��4`�����~��KH�z��P�Z��҅!���O�%����z[XQ��|)������K�ۄ�4�:�7B1x���o��>�6Gn���DwM�u5Ū��G��y��NК����j�9#Ki@6���k�(�.,�N�yS�K��CGH7�����=h�BӪ�0���hP������8���~�>%3�\hp�Y�w
�gDB��Ӕ<К�)���Oh�&��3��� ��7VK�/�ب�Ǔܴn,H�rR~��>qaj*�"Z�-c�����OMIn�h��CgۢAj�.}�.�E�)/��$��NvB���7��@%�y����WR&ۜBC��4�C��|����JDC� �Ѫ>�}�����F���"�o4����4��I�!��W6�E����,0�Dfz�N{�O������}���9���!%�&_Ĥ�
i�ψ$���.�n&昋;��n̲�tt��uT$8�d�x�F��a�$ix��s����X����o��/d���{��zrM��Dw�fl*VO�۽��rޱ��V!P$�R�MOQ���c(C��C��HZ���l9�z������Tm���Q"R�Q�N^, H���A�S�b���]`/��n��_\m
l��٢Q�/�p�T>�S�]�Tf|�lj�>	X]�Z؇�eD
s��$m�����	������&P����"ûI�(h��k_|�Gq���wZtDY>B;�B	o�D~���2�l&���W:�¶ی{����sq57U��+agf��c^db��4���Wm��S���	l����0tVpGxLM���4�YgD��1}�Np���F��Ə����r1+v�mԞ�p�x����_������F>~���W�'0�L����+b�ZL$�������v�=j%�a������92��>�M�	S`�ХT�"��<QB�����%�K҄p������+����+�>�!m���D��\�W"�Gk#�!�D'm�{��s	e\2;	c.vϫ�i����iոO�t5\\x��w��>��Фz���%6A����۵1���<���%}�辆�@�-V�8ɉH�P}�ɯ>����S4A��X�}�V�TwꣃҦ��Z�+�6���x�^�^�ԅ���Q
\�A��I�88|�yV0�T~���T߻�>�m��c�&�X����J�]��@���<7�l�]��Py�XXskii	X�{�F��W���7{�� �����1j�s}������U)�A(�
�����)/1әPq����@ⴒx��p9�!�����Ѷ��K��c?�{�-w�?unԝ$MDI�ô��z õ�G���Il����R �S���l�ZlєT�T%�^�X+�V���L�c5�cz�)TGh/��;�P%���.�Xh情ع����.)�G���n ���:�,�_ơ�OH�9G1���kc�pU�{&�j�̼B�lU��J!:Xr�ig�qM`�����&5�n���0��)�
�D����\.�HU�L��O{�'����"�jV'=7�v_D�I��U�>��5�,�#��3r'Y=H ����W�1Ӌ�}:G1�6�kb�H(3PGH��gD`����a#ju�����J����2_5���8�VB���F��b�܊�d�G멖��#P��亾~�6ja��(���iA�yz>��0���脮�Kui�^����� �d��jUs����޴�+՗�sQ������fQA<R�	QI�&��/��2����f���Q�Q����c��{���s�،��
.��c��4��wj�#���i��HG�)?��j�8�4�
fj���Y��N#�5�U{eq�é�UhY�*��HOfU8G��$d�9���?\ˋ���X�M��`����wAכ�缈NL�ڐH_ ;8��)~z��Az������s'�����=q�{Z��2o�Fl���Y�gQ���R���J�Y��t��:�NB�Mh6%�����8d>"3��UQ�м����y����C����,Tu``�]U�l_n5��L��Ѯ�Œ��-��f:ܹF�pH��,�n�� �f�o�}"a8��m?�>�H��DU�eFa�rbKgQ5��*�٥������UHük�>���5K�٥���˦A��sh.�ܘ*�Y�>L)�h�'�q�7V��T(��uF��m��r��A��ʰv�����������U��N���q�<�lk�
.��?f��Ν&��t�$\�ֶ�����JF-#��5٢�{v���_�?�n�`�IJzJ /)�t��}�Z4��3��GD��	�s�� JK���Xeֵ_S���"uo#�Mb�MB�r�X�*����M��wf�vK�I�]w�/��|K+����f]|������X5}訅�)r��ڀ���1�[�k~�]:)={��$kU8�,�e����˫���ҸL��B�ܻp�
�EN��F�l��t�A�� �ٴ2�U,��d�.����ug�g��;�nR��}U���#�A���Ѯ�1��	�⮈l*��Q/���r�;,?��Mn��Ť&�zih-]QK�[���[ ��� ��3��bB�o�m:��Ґ��� ��SId���V
KG�&�s�zA����D����u�7�3�7�K%��nD����"��% �[�r}��>�*@�������=g��˗��"�����Q����݄�	{��]�m���5d�S�{��OGUg�.l��ODܤ�=l��E>�� ���)�,Y|R�[�45��Bp���+{��7��_x����^�hj�2�A!:��uR ~�m�#/�v����^+?Ƚ�y��Q���:�1��<{k��\]K��9�L�L�U�}�v��9����sv�~Bm��2UR&ֵ�*yt�R[S�W��ϒ���C�>e�1ldfq����ou����*/J��נ�z���e�ⷊ4_/\!v�+�&.���L�=-7íCV�k>_<n��wMg$B\�`�c�����)e�v��N�Q��0��^�T����Ѫl�*Wk3�;��U<�˳�9�\,ـ�I=^1�Ƈ�׍�jO�KKn+�6[N�2P�f�&�=��XU����_��;����L��d�G����� �%���R�c9��s�Kc����x)V(���W��E�\U#�-{~?e*��*Y�=_D���F�����pn��L28��i׾��C̨T3���ڎ����m�L�+�M�/S��y��sE�Z�F��A�(��s~��?�'v������I��1{]�~~��S��+��t&8����q�l[��S�h�� ���3^X;�(���^�f��t�9�v٬�}n��Ô�[Ted�m���=� |���I-K�B�8���;�
Y��G�Xˡ�	
����}�w�p�_��9= �k��%�n)"Y֋	x��Ԍ8�b��Z�s**��i ���0�ب�w\��$1z�t���=śɨ;[}�O��Z9T3��6ҁ��_�V�[:�_JU�	lVʗ�.`0_ok�1k�n4z�[��ӚH���ʋ]�X��QA����Y:����#+��pP���v��,`���*b�'����ۡ�}T��N��w��D$#��i7iE5���+�xb�F�����`�u. _�
��^������)w�S'��L���J{�*��#���|@��x��f9^���;ȓ{�!<h
ʻ���Yα]�����)�2)��~a"���&ݴ�J��w��^��㫵,�����Ȭg��<ct�d.�+�I/���pd��vc���J�(ע��1�K������fς2\���- ���h���� ���&Zt�
^��1�xc�v[{�H?/��<a.�]F<��;�k��e�Hq��NPv7\*������X�o�*���Cף��/�O�u���H1p�-�ȕ*s���\��	���>�~#��n<���;�p:za*9�-��/u�Q�(d�p�N��[X����r�)u&÷}�-Qd��5q�t��gnaO�n��Hž�Лhpv}��j	l��E*ӻC߫������L��� °��Z�-�:���X��K{�����VH�Ic�:�>�=��{����A�������N)'(%����XJiccs�:S�<"�����a���$H��K���<
��!a��A���!�:2��\Ň�����-Ee�xs�f����~�!d΃E�>^�GO����[JƤ_���q]����_����M.2k'�r� ���pBh�z%j�l��Yk����M�{h��W-C7�{(2��:}(T�=�A֯B��:d�~�U}GȸY{@>�N6��F^I�L����VJ������rZ�e���)��H��)$��(i�C�#��]b�ٳ��},[���E�( �R?�,B>��h�N�� x����)�d���#ܑ�����beAB��al�D�m�t��(��(������4Ƌ�U�Y&��u��Z�phߏ��櫖:|�0{��s'������j���φ�������VU4��=���aS��]cv��� #�J�Z���T�)�8;��~�@V�
��v��&r��oQ�}�~[(x��I��m���}*���~EI�PZ�B��|ٖ���$Ձ��xVǱ��/$�bט�ya��	��ӛ`Ѯ9@��޾�7>>��Yzhv�
Vۆ��x�)�kna~僇�Ё����Ď�}z������3�6�]ת(bEN�Of$����V�����
sCV-�'z�������A�i�60��� ����ξ�^�[T7�5䕙��\$ٵ<�ӵ�!*�ZaҴCD��;+|Xؒ���O�F���a�ۋ��g�+f�U����]<�<@>~xn�/����AW	���A@Q��k|�	�Y���HD'V�--UÞ+������+ [Rr����|��<�S���W;@����/�Y�w��WT�N�����eO����7�W�q��fCC��������-Л"q�k������� ��N��+i:�� 
 ���P�R�7� e9�l;������Q��i��V�"�ت�	�I�:^ZWH=�pfkZ�⅌�V�d��<A.������_����:��L�j����I��zVZ
�拴Bx�+�{�ϐ�7C~��;���x��wz2�\?��8��X��(ܘ�|��̨�4�ɟ�J����˘�Eu M��H��a�k�����w�'�܅��q��\�Vc"0�A�����k�g���)�l*��/�PyP揊e�~�Z��D�}��i�y�������9��~���{��~�D�G���Q�����m�a��*j0\�3���wχ�le?4��S��������&�0�˭o�4z���v��l��yx���#��#I/lL9����]e�V׌d��R����n.[��Sؕ*N.Q:u]YI� ������->��j>�N-[n/S^��n~�WS�:��Z5���bf���f����/�);&��IV�����u)Ҵ���}�g\컰[I�l�@
����<��_b1��%vv��+���`��J�c��Ĥ��fC0�;��ގ���
WP�����ӵ���s{B��q=�/5��<+'���'����w��l�b�ڑfթ�$�:۸'O ���{y�h����9��� |w�M�E�'�&�:��ǹ}E�'�˛�t�̩I��Y���o�{7�ST��J���`́2{�^!��?Q{39�d����BHeߞj/,�U;��0�g%�^b��B��9��T)�u�2�B^�g��F�G>le�O��:����	24�lg����nͯ��������%a�ƌ��G|^|���}�'�N��|lP��{Q����(�$Z�\��9 ���i�_������NEz�F[���ڽBo?��Q��ڴ�B���� �yl1��o7�<�F�a������	M���eѠ߽w�|�- y��-�K_1 	�ZQr��JV(�z^��![{� ���A7��n��xl�:L)����L�� �IeUY aU� �f��i���4���ѳD��{=�X�������*�;4�8h`�d��F�xEQ�tB[C��W"2V�R-^��<�����'���pCY6,P�)m��WZZ �*����g��|�������0Tn�j���"�>�A�g�F�c7嗙ܱ��S'��xbu�X��hk�'V}GY��}V��9�ff;����]l��V5*�s��׵;��ؤ��df�?u��ri�$$��r+�*��:li1<�ʪ���g����ڵC���4�����+�uodd�5��oF���4Muc�A:5��I-�N&G�`���`���7�v!aŖc�">56J�]�t\�"pо��5�>�����ZV��:g�#��Z��k���[��i�Q̀����i~Jk��>�E�T-c�藠�B;*����厨��f ⺼'/����u�r�����G,xdV�~L�E��>&\|�^МJ�|��5,/�{��L��"�JC5�xq��yU5������bW����\��*q�1DH�riJ	��~ }����;[�7�)�1k�ʷ��iُI�C�P--���j��e���{�Bl�Z���mX�.����N�������#U�iK�Icv"�+v�\,��/�O��܋ϐ�3q-T��U�/����$�ȵ�x�tAiFN[A�S�!K_6�4Jd�0�D!Hȭ6!�������Ʈ䩾\���#)Q���%��8ڛ�=!� H��+����9V�.o��dV�`f[�ƫ����ѧ~�ѐ������iznn)�k/���ǧ��qEf�)l[{6}6���+�,3�l9V�U�����0J��Z��<��c��E�J�(r P`n�W��V^+ EzP�J�=�!q�h���z�i���壴|�GݮQF���x{��:�u>ɏ "�ɪQ2�!���:s��S��7��� Ȑ~�<�o�X⫏�:iik�JUR2���	iX�����x6}�ߧy��?8ݷ���5����ҎR5�P��<��P��(��uD6�ߕ60H�F���JJT�5q�m�;�8�
��5�GO��g�ǎ�3`�,�o�����_�E;��+�xa�R��xD�v����7�rNNN��n(4�L0f:B����v�#W}p�Z@��6�����n	�K�W�9��*\_(T�'_��u	��Hx"o�{U[�̝=0���`c�;���
���	��@��!��������+�V@�D�Q�<M����g�jE�!��1�};�VZ��ɬ���qo��k�@���T1Z�hi'�Y����gn�ѕ����^���?_x�e(B�<+@��W��-���,_k�B�)�gef�$��5���?gH�'��1�����T��|�t�bl�m�q;�[���C(�rR�o��1�v�zz�U���Ha��#�A8^k/���VV�	E�q�.�̙/99�O�&.��M[ tB�����������@Wg$�z�#�eo�`l����kN�񐡛D�>m<��������Q.b4Z��\l�D��.�dFTdE J�(y�Hȳ��e�˞����;�ڶ�>������/��a!�o�m��^A�DK�Sr�	h��xU�C[�&;_�Lv@�^���$\���5������U�})������mH��č)7���r���g���A��S�B�-����U&��`vu-�ޟ��b��GZ:���������#��D-(�-�Ӹ)���UF��.ZQ�֙�9��<{��tm�y۳��sL�Dq�uQp0;��tEG��r��k�g�yT�ٲ�T�O���}��DI��n���:xh��M��j�}w=�cA* l �9�����D���q���^P%ۭk�� 0+k��o��j��3���#Ϣ�zb��r<] �+��U	&�����%����EQ���k�`K�g����t��0�<��-&���Y�7��̙��硻��%`I�0H<-�<ip`�����N�v���$����>E�b@���㆔9�������k		<�zpش=���
���o!��|�S�������ed�$׉Vm�F�Eէ0���,���ll�Q-[V>ā��{�&������V��0�/�q���dHf����NѦ��źVA[��x8�̝	q+N� ��J⩈�m.��dz�T�X�\�:���������#���]�ݎf� ̖�s[�~X���J	�T�bQƖ	��m��$v��������8ъ�U5���P˒g�+��sx7`�a�-Cj>��տ�W�d��V�5k�j��Ӛ�0wP�#��+��o��ڊv����.J �S�:��jV!�$��Qm���ů��)���<�c�#��V�d{�o܍�&2�P�,����N�~���b�OT��
��1Ȕ|�����WDejt���5�fj�Tm%���=>T���@ς�K�qPXʄ���}������C�\�`����f��ٕ��s	25�=r��J��� B&7�K��pzS��}%0�*��~�甼�J��Z$/Q�"W ����{W*�S���QBsͳ� �C�X��r�"R\�}�WX�����-�����fi�@���[@R-��$bLC8jbc� bz���{��|�ѵ���ZW`''�/��Ϭ��:3���߼&���!4����q��������Z����\�Cy�iҺ��"��~Wq�7�Q*�v�^:s�&��ٽC8��� �x�	�����^��BS��3�R�!�~��gN�lm�|q-�3�<
xo��b��:8�L�?�r��F�S�����MC����fS�yr<��8{��������Gv~ٟ�O.K�x�KOd+�' ��f��E������'��K��<{�oIk�4����5���]cQR��1�l�.OٽcYa���)�Y� ��2����5��(��3���z:5�dH�w��NA��'��. ��O�(�HW2�C�YN���)���hwn皨�*�yO�X-x�>�m�~â��Υo!�r�э�����7��5�NOIp���O�K�CLw`]�vmD�>�vc�a��(; �u�-c�Ue�{|�=�9A2�c	��^��c�G���ִy��{���0���s��56{����dٓ��eKH�)���v`����[�Y}�Un9q`��oA\�}����ـ*��`{�n�r
ٴ)�.r�jc�Io5�/��S�F����;�����(x�D�k�`O�OƖ?���YQ�%4s���J�զzQ�[���E%x�����a#�qK�S)�}��D��E����ڋ�3W���a���*yp{�eF�,�}k���'\�PG��-���W�'g�8'�F�>װiv|�t��2Q5�g2.��ŗI�C�ac*]���5�X^W8��)��#�?�y
�<�~��ss-[e�+:XZ�=-S��l�:�6�sc�{
}.T�8��%Έ6�����T����?jW�ib�;�&9U���7�GEy(�TcN"mq��
ep�1�  �'�J�~���3��8����؏�P���Z��:=]ܪ
%DFDs��}��������%R~�cx�Mp�y�n��ǜ� �QI53墵�4~��`(���n$�٪��S+�Cޒ	��>�ՙ�`����Y^)YY��N���ݬ1^�l�̅�>1B��Dcι�x�\q��̍~Dz�W�P�.B���uWU���b���_�H{��IQ�Q�d���c,kңW)8�:�6�-�P*��7'd��eq��
�s�I�7���+.�G�,��"pl|�D���p�6�76m���������9���_�&Z��̉��{��K�	��P^K��SV���߄�8�Ȍ�Z�Y\�NG�Țg���Vz:5�+��
���K0�z���r�C�����4}Γ�g|�(�9���aɰ��i�M7xP;�����p�`��k@M���)���߮�7ݴFKsy	�KnZK�b0�e��tY��d�%KaA�$yũR
�CMN���KBF�����bh�>桨��q͒_���pL��/�h]��|��
�,�1m���7�2�~ $�xDsBS��݆�=�pS @�/����i� �h�Y]��ԗ���� �o�bŲ���D�l����@��G6օ��N���xHD�gc``���������z�#����Gcү+�$'�B��"�K��5ޘ���K��R���
�Y��mU��
f��ēc��q_�݁-V�k�$�)1IL+�Þ�B��:�lE�Բ���_l��Փ�$�,����x�s08��vl;�ÙU2 �MPz�Qi��>m���p��?+B�g��$z��c��\hІA������B�R�t����ޙnz����B7�|���e�U\L�X�֝㑷��:������p̠|�s�3h���^��K�`Z��? "I�܀sacJ,�iu����Z�00�L�}-!��{���
52N��t�;/������4���B^���r�A��.�i�*��1)_�j8��o��x��V]n����EƊf�$�x����A!�!�����x��f:�@'r���U~��6��n���ݽR<�����S����T����H`�m|3M���GJ�LĬ�/��ZH�+|LQ�b�~�k�D�0:n����T0m3b�~�(��.��qj7:�v�#�� ��,	�0�n|�x̙�u����������L��c@�Q\x.V|$R3*�x�#%�����k�U�KnϷ�Y����~x�ΛRa��� ���3[����eN��cf���w5y�H�����8��`au��Q7~y�-xW(�Q(��U��"�ǜ1%���WK	���+�o�R1#����
�J;�WB�(y'h��x�w�ֳ�o)�p���ܼ]�I��C=����D�4�̑wiI�V���,�(f�t��0\�[��-��
6q��P-��~E�{�g�A��_uCY�ٴW�cQ��̿�Ʋ��꜑��J�AM���7�~�w������#${r\�kS�.���m��@�z0�յ��� ""�?��h���$����~{_���K�������yU���f�s�{�:������K�z�ͱ�UVǫ�S��0��$�|�Y>EYB����G�6�ViF\�>G3�茣��c3�|/a�_�S��1|]�'�F��T�v�	�ý,x5�-��r]T����j2��J���W}���+΅�m,v6K1��j7��?��Y�E�fdH����f�֤no��[��9���f��ۚ�x��˧��9�d!^���.a���nvC��~�e�{i�����8_L~���z����}�喠�I�1������>̌W��7�UM�/�,����� 
��M7!���
+n#)�p��.�}��H�U���+�	z	Vm=d�2�>be''gD��Co3՞��P����y��P��_Z�@q��m]�8x�������v�"�پ��j/�nY�����
�j�1�^�1�7?tP��Θaܒ|�������Kqg��~�Ť����7f+k��-�x���
b�7�������,�g�1d� /_Fh�]*7�w�'������m2�f9���YZ��ʝ&��bH.��{���O�L�R%�5e[��c4t>~~�:9��m�Jz����d�n&��(f��2f��������2�z^]�F�93g��K���a��H�4]���W&QUҮ-��M���D�v����7//�����w���C��\~���,L�[��{(�Õ�C\���֫9��a{�r�#�2U+g��/	��I�&��xL�	 YMg?�Ҭ�?#�U��)��A��h���q男P,�&�e���
�5��@����јa�J�볷�?;5kao��N��]�sN�E]�G�V BI���")� �RM,��E�})H\bƆx�N���9?�́oz��֗���~�ݩ#��Xո#���pm�W���n?r�@�֧�q��}н�C�$����-M�P����1A�������7U:��#�ŉ%�|�F���2�_,�Eo�Hz���4�Q`)���KR�܇1a5��������
ֲ�΀�(�m��~	��B�W�.���{<W���z2���h�I%�Ȅ��+2"�~��d^wk�zT�*�U�v���X�j��ڑE"HI�}qzؾ3��Lڛ}�.>y�v1߇m�`T%iMlv�B�x�u�7k�T竴~���o��
L(<�<��+e�Ǎ�7@����Nr�r|��̧�㷸�}��'�r̸�}�*���^�o����Lw:Iyv���Ƶ���w��^����e���^���CȮJ0�|��!���}
<�zI/m�E	�����3�i*v��nŝB�	Ǣ�`�$����oZD������k/N��C,r�O����Q�|�v��rPT2?/�7�ji��@�ALb!N��C	gD�xh�Pe��f��kk/��ػ���3�D�,�t�й����ý�OAO9��#w�#�<Ρ��O��ǉ���ͻ�G?�<Kx�0hn)����|̾銉���NH�?���e�G��ΘD֥���Ău�;�d��2� �*ȩ����Ky
S����^ί�=�̵�̎�_�B`����+m=QK+�i��>�X�������3�M��?Oj�%���VM/�$Y���I�����ETX��e��{#	�B�W���~�"s8.�>I�e�{��t���`�RY4��j-��#>�Yմ�wn�;Q��b���^x�z���"�r��&@f�Q�J�3�ه*Â�c�i��v���ޙ5V����~F�<�9Nf)�;Ҫ΄�4�H˞�� �WSB��E�ܩ���.�[�T�	���I|�xy֬Dm{YW�ݒ�]�ٹ�Ū|M�1�<knkS����<M��Tx��#`Y��l�>i!S g�6F˿��>X��?��8 v�w9�{@�[�_�T�Q��h���0�ը���ߚֆ�+�Ţ�e����.���%Z��va�&����浌���U�w�=w`�	�Z�^�1�uSR��!5�<�#S��۞-2�ߠi� ��B*���s��stf2�4��_��KN�ڻ�b�sN礃���J��">��}�[;u��?�u��T����^�T~��l����nI���/�o����ϷiW�Y~9���,�K�ȹ�{����鵸�@4šȷ��k���ݓ������ŗ��
��a@��7uo.Tiɺn�.�cW2QR=\k5(�1ef}>ѱ���+���ٹ���.{����1��`�c �ߕ�a�S(���_�PQ��m���g�:H��!K�Y�66�����N�	o@^晢�'i�O[��-~�^�B��a��삶iAP�QD���A�����WQZ)i�X��A���A���%�{��}?�z~�p�sf���f�9������IUEt�Ml:Y�W�6�E�h�y����ًF��$_�V��
BA9��G��\�s3UǊ�b�o��E*�g�3=�g0iթ.PD9��=���"]]��7]�<�̙��<j��.���6ƶ�����}\�'4����lԡ1U;e,[3��y�S�Ə��p�tQ~�  )������I�
��Ćt�@LM�����G�w�3U�4O����>�L��{�*�:��qH�A.Nk�kS*�Ur��U��4Tq~$g��,X�'1)���	=���dG,��R����Kp��ԄJ�*���tQ�;�bQ�Au}�<��PR�tj�Fe �J�"X$_�;�Dq_F��< 
Es�d� 
#2�o<fd(������ؑG� $eg����I,�,��W#�O!F�[Sa���8����_��U���p*�����y���,���[������
�	�^��{�A�R�m$Y�ٰ��C�-�э��c}�λ����IϷ{��M�'FKm��A�T#�Fʖ��zZ�<��q�T �sS0y�A�z}���ͣǩ�=r�ԁ,���,��%������>�ʌҳ�<G|��o�	�Q�]���΃;3�O�]UF{L�&S�4
�Z2�r��T#�{D�L��W��Tw��9������ȓ�Z�c
�ؔ�
}D�I@��z]���k��hk��Z����*"��U����P�R1O�`�C׶�h����{CZm��J.�zE���ۣ��Y��3����X��C�����vF�p�[�5�[�|,��(cE�ḭ�ߗDio�����1�R���0~�Vu�A����Vُq��=�a�#gfNue$]��;�(�v�~���C쳵Y��R�$ �V���m���m��ɒ�T��?ʏJ���QWG���p����$k�L����b[���;�!��V��x���J��٘hk�����1�`��ͺ��l�m�=[��&�Y�^E�bfwא�q���T������������s��̡.C�V��x�)�<<�x���L�q]B�`��z�W����1w���-������������.��Ż5�zH��;$5L�ފ�I|�/��뤱��o�ð�HOZ8mS��_sG⇖	��\���M������r9c���jA�D>��{'$����Jţ�>n�ly�?1/Uz#0F�)�^IfU)~����n)��cp<TG�������ϕ���b[�k���ht�)S��J�A���{>~��A4�T�ֻ��_�y�5���>Y[Ðw���M���d���>��ι���:k��#���?<���>���0;�3����m���k���?�dCr��"R�o�1�Z1��v׸��@���^^���b�=ӗIO����m�J^Q���o�t�r����{�,�0�߼��?�T�z� �H�+R=�L~��������6�fo�|ڼ)���N렅�%[��R���Q���4��sj�Oz��ڸg�@:�AF��x�n��Y�X\6�b�)]��0;J}�[�����g!^E�Ӥ�J�)�'�@Բn������Kկ�j�|�޾���;����C*�cm�I��)o(�^S4TZ>d���g���S~�<Y�m��l:�\�y��FEm�*�<}M��Sw`*��lޠ�I4�#�^>%1����^W��8K cz��@/=�b���4�z�M�2A׈M������j��yq���-/���$�~�d��UV�3����Lbo�S}��:.����Ry�^����E.��Wb���5���>-����m����� �5����<6���xH[�4E���&p�ܼ�+������pJ�˱6�M��Z��;4�t�lX�����o}C�d\w�f 厅Z �J5�ڂ�������۰㳵�sH��ᇕ�|rv����܄K���w�o\��B��G�YI�x�`B��F��	1������m���ͮ�H�#�\�g������=��]�t��ɚ+V��\�r~Y�ݍ�VA��	��-SV/�e�Y�5�p�UHN�)�p�^;j�����N�%&y�6��&�{.�Gy`0��w4T�$6u�ʹ�F���^nVұ�KCy����6�d���h%0zK�ͦ&��4W�"q����WX���Fɏ�Er�����8=�����zմJ*�W8��`!b:����ٯ�z$8<c��c�Wu����I�F���9EE���[�ۘ^��N5��Y&��y�>����2wO��Be=���pU��A�1v�y9˽�G��݀���_��%IF��{jE�������kqaZc���c�i,�"��1s3Z��`N��\��D�{�Ƣ<y���?�ޞ�5:����+�+������Wn�I�e���l���hC�b/�`5�پ�z>c�,%�{��W�=�˴��+᧠�&n�r���)�- �8x�0�����N�[B��]j0�o�P4�^��h^B^WV*�^`3� ���vJ�7�ϵ�}kdEj�h1vW��D���{�u���"��Bʌ;�!��O��A�P�uf񗚜CM:��N>Y�Ψ���,�J����W�13M����_�]I;pp�,�|,{����Z�+�V�c�aV�� �����rS�܊r��$�]�!^`i���c��Es�*�?��Q�����z��IQ7;`�gz��cё�`Qz�v�0d������ϑ�]��c��@��\T�*���m��.4zjvZڋ��h����g��<����B������/@S*߱^��sY��>��d�oʝ�}��V ��s�Jɯ��9��g�^�����n�'3x����	�GFr��P\lU�Ɠ���@���O������b���N���A��ab������!ڣ�g�ݸ����E>�΄�m.����?�Q�p^QC�w`;K�0����\gc�~X}��D����mre�t$�����Fc�˱O1�V��s����E��Ru�hn���i���Q�^�$$��a�|X4�����Ý=i̩��������nߛ�Ol���QȖ�,�M����Jl��3��������y99O�J�R�~�1��.|��R���]���Z�Zn=�}�v��Y�!++[�����jY7������t���a�"�l�w""<v�W]j��1�����8з�-3��̯�$~�����wQQQ�{���ë�e����Մ 
66�xn��L6ଇ��uL�Ė�o:lO�P�^.K���a�^TL����Zݢ�j���f+��w%��`�!8t��6\`K��R�ô�S��u��gn��is�ؽ��8=�U����c��������ϡf�&8�r�aY	6}�7(%t��NWX' S���""��=�>U3Mv�204l�]oa�.��
J���3@q.Ou)f5�~(�Gu��ø�viׯ�Ѷr����S�<PњSv���vq/���»�B�0���˨�	���	zzz.X|<��� �Gq;﵉*��߿U\\*�=_�|���p]_!��"L�#�Ig�F�@�X�}|+p����q�����Џ۲Gyi���.n�()=D9�������$��AV�#�M�P�	i�{���'K����1�}�S���Q�Ĉ�>�"!���aμ��B!��[�f�k��Iͪҩ2�?{���_Ĉ��e)����)H��r�Q�?�,�Ĳ%��,�l��;sM�Q�$��]*9+h�-�u�@�9Ѫ-R
��qK��C�rA��P��(�_���O+�:(�y[р;��!��>
Y�ߣ�
-���)Ay�$v6�l�v�#o��f��3+�x<�8+5ǔ�Z�k��}yA&˱���X�$��jb��F�E'��o^n�ۊ�$��!�$W�4ď�_�	nwt����=�14�b-�Q<�g�Jg���-�QE=��SC}������n{��n�{�)L�W��X߹���b��S��l�3߲��ы_�XǷ���9��1ԕ���$�pw���MpH6�=ju��=L7� �2�x���t�s3��mPZϷ�3��Y�Tt�S/�V3���VD@�
u``�I.�B\z�[04����[+e�~1t:K ��'t��5"�k~=�;�
�dLܽ�iyV��t���5�E�j�n.�K[�B,�,u���ʡe$��T]�����i�vE����=���s��1��+.�7���[ԁ��fl@�l0|��l~t&.`q1����̼��A*�_��[���ٙ�+Q��짺�LE�fy����|����ۑ��J?�l�"�����|�?��@; @�*�e�����Hr*��+�Jč�xx/��쬅�Hh�p/\��d1�����bq��m�.�w���t�u����5#����k�굚�9���sa�
�e���G_Kh�U�\�K���\��jN�L	|֑�P~퀍���� .��W:nFa��~B-���;�b`��	����1^��Ǔt�t?�a VUzK�}|����hVpx{ﬡ���ao՘ֲ��a����^� P�qz������),��q��W�݋������,IY`�;�)�4ƵB�^�0J������\�
� ٨�L��Y��;]������P��Z�Rގ�g
�Q�M�⑵e*"��શA��J�o��7��?��Z_�F�*Sy�)�C���<�N~�kT�v�˵�S��/�V<��R	K�o�bӰ�N�?�i�<�۹�H�{l�
�JLˣ�p>S����*�6/�.�O��g����o�'��6į����m��P�@RAun�DIZ���k,=�W����O թ_����L�IQU�k<F�j��"Ά�@�;��1ud�z�@^�#Mp�;)9[��Bj��SC���tn�Hu�0R8P0�l�����E����Yii����'�{F�|�/�v�P����R$��6��xb��Ly�����D�l�GhZ�E�u��;�>�iE$_C`]K��P�%9p@&?�^ιq���_�~�ӡXd8�D�akь��1-�1"6s(6�gaEHP2��uO~������� �\��"�^�ۊ��-�ޖ�u�r̓�2�gUp�q�;9ux[&��B��0VÄi����~ͤ)��'h��$�)�	�+ۏp;ٚ��+G�����J�H�wUXI/0�@�rt�,rT1���}�|vN-EDd:Y'��:1�4p5)?[(��iS����K�8���䰰Y[����^�&Y�~x,��	8s���%ҫ$qp��cczH?�,��f�-��K���'$�/��9r��y��s�i�)��҇L�[S!�vm9F�#���,��g>�/�.��z����H��D6�ax�۪:��Ȧ6*B����o���z�_`�q#%��;I�K�%�g�_bu'«���OhH{������{����OOX�Z:�j��	��|[���~�1gk��qD/����i�؁yz��@_�~q�2퟼�NG{�+�����}&Y؀����1/����^0KU�V�Y����=ju�ޟ�RȰ�j���Ϙs���Z{F,��SI\;��g.���O��`�y\����J/ʓOs��.iI4��6����?L��E�怇)�?��T#��,}`�&�+|X8F��>z
GK�<�K�}g2���h^�VJ�Jm��M,p	ûYw��u¾>5~�j����C���$�Bg��Q�H���v{Ɖ�/�7�5��M�,�$[�Q!��R! ��dqPD �Kv�[N-��r�W>�y���SZ #�jˊ��m����'�4+�ǧ��k�>�4"%T���M ���o��(hݗKƼ)�E�t3a�%�,�8��Y��Ow֞�Fmw;�=^z�a*�h]ZJ�Iɷewe)��'6��m\`������adz�UǴ^Êצ3���.�K��G�;Lʐ$RRҼ�B5Y�P�k
�R�oi�:4?�̱���Q�i+��6� 㼔܏3�C�ɩ��p����(�qśO�Y�n��(��m�	tħ�ho�����<�(���n2�׆(ǳ��8a����u!�޺����n�bܦ?�^��;axe0����dw�����4�J!���Ha��6a�c�*���h�ؖ��-X*&�ɠ��u4U�g.-b�c�s�>���[�{V��|����ݱ����ITB��d)��O��D^�۷o��&�<�����mF�O�'��\�[p?��r-:*꺆]���`�6l�o� jߞ�pi�[j%���I�~"j�SSQ�0���&1=�Y"8����Z�3�����K4T�n�i��.�@���r�Qf��!g������>[�mrUuu\Aӱr�&��o���ԫ����]���[��_s��K��O&t��x�h��5��a�7���ò��N>�U["���e��_o<��P�yM������0e�,�e[j�s�7a�ԽV*�;O|rn���>G�u���R)}��5KG]���V��#�v�|�!�kf��2*kZ@��V�OAFe[�f�޵���[���l�_�֥�V�ą��(f��)�"_�;���D��p�
$}�\E�N������{������}1�5����ëO�V��~=���BK��h?v�.R�ר����ވq�|k������Dm�/���7`��c(����>�
��p��d��^�OϬ&� =���ċ��w'6D�h)�M��Y�O@L޼�!��.�_�UVΒY�;HL���yɷ��cޡʿ�2�A��5�PƟ�Je��RA�j�[≂��ؘ�����W�SZ�$UI9]�dL�~q��VS������	����>�"�>���l`�Ԛ������w7�zt=�s�ȹenP:E3i��S]ӕ��($)�N�C'bA�XA��uZ�b��
������@�_\>�\�a�E�QW��'T�*�xa�9-) ���OLf[C)x�|O�S���i[;::_\3.�D
�XږǶ���Nz&_v;B0&�(��
����=�+d���$Ȅhb	�L/j��_0p�Ν���˟!~�F�6�E�G�Wow�QSO���˓��e��>�\=�(���j��ʈ���n;�5�����x�EUm��6�{�0���� ����w;�����ϝ�.ø=��a��xe]
���q�k���}�%4;.Ƿ�hҮ�v�x��}ˀ�ΰ�Ԡ+��j�iGH[n�z�MiZuO!�ڒ���cF��#V)*O�Jַ�JzV'���{�]j��rMX���/��ws��OR�����'>����й�������%�?Ed;��C�Ȋ�)4!���]��c7��zIW�^tcC��;��te�}�<K�ɱ��y<���9���5��I۟/�d~xx�q�ي��ݢ������G��x��j��A��0���m���7a�[� �j�����!�=-\:t�R���*9i����(K̚��ȴ	l��j����f�_��h�O'E����:Z�P]`��C��!] e�WU��?��P��"o�+	�9׺߾y��`ҝ\ ���s��j��Iz��+� �a�eH���k��%�=���צ.5���⯠Rnc��ep�jZ)��M9�ݢ����[�0�+�F�Ry�ש���������5�hk��m��8��ݑ-TTT,�o�.$��������Zqώ����X���70�z�K�;S?E�շ�!ݮ���>ۂ�a۰�F�g�/..�7D�"R^(������g��g9���E����z�w���Ҧwm�6�!+a����ǩ6�;���n��񱱵�����c�rm�h�!�?��*f�;���k.��Bl��ӻ���XH�/��̜?�t�iW���99O;����֛�>���|��칦��o���˙��a��W^@Q����Ra��ӫQ��81���.A�ED�b�}��q���q���J���z )݈$��YZ{.���.�S��K��m8�?�JA'1	���u�[d��*�|�����5LڬC�6��8��>{��J#�|4�)/�̖+���4��l�c�6���8x	a���� ػ�3��Q��,����P[�P1������xf��g7o��9����&��́/)�ߵ�0����?s�|�]���,n{퍚V�����"�\�����v��NKŽ�I��4M���进�)6�5s�����NZsD0>��T�%�1��gx���>���Vl�>znn��!X�D�����q��JQ�.�魢d��jgdo�������Wۑ�?��IT&Jqu���K#�Mҷ;,U��۞�0vbutk�<��4��rW�r;vhq�a��(^�LP�����n4�'<���zP�l���ޠ(�5���]l<��U��{�&�N�b�k���[�B=��h�'�V�.V-�3��vꩱ��)���mZ��D��-����*�#�,��m����)g�z���|��N��sv�ݙ���>�y$��Km�[������3�H^:iwbtG�*�1�t&���z�����	y<2��� �E��Q}Yop��	�L�窪q8_��m���������M�v�666�ұ!zN�by9��+��OYǨ��t��c��;���a���	���T�3�~OL�9�3��a�`=>�B�ciNңL�fhApb�w^8��	^PP0V3Z@>Q?6Mr�A6g:�^dT��kD�^�GDEE��k&M�� Qř��s;�td��X&0��~�Mrr8e4U�5Z=�9�;"!n�Bo�s�Ȋ@�I_���/ ��Z������B&\VWW�xS:��2cu�՞*%�/��sYƤ��U�O9"-���cK�J�^d�"rKk��­C/g����l��-�o�l��T��ļ�e��{t��Y=pW��C ��]��s^= \�����51����Q@���gl.�jyŮF�����]��iJ�����$�����*�E�N����3+����+.�U���[dc#d��_�:<&�I���r`��>��oVlM�ȼkZR�G��pS�z-と:��Q�W��{pʡ�+{��m�ψ�˸S����-�Î���4K�+d;c1�W���i�����k5Χ����Dt�h��7��Y�)SOk�F�~G��)�E�K�+Z�0_����l36�����}d����α~YfŌ���[g�a�z�6#�CQ�m������v���h�NT���P$$c7�&�7��{v�9�<�c��:J�4��p���N��|�����Hq�M)J"��Nv�0˂M���,�)�x򇕩�~���ܽ���t��j��͠�0A��ix�>����""�������Cʯߢ���R��8V'���&��p���n��!<�B��U��v''��7��p�M�,t&d�R��A�Y\L�g;%��I�lJ"�Έ�l�O ���N'Hi�G��C��g9 ݡJF�Xďc��|ׅ3�e�z�71pU��	א�pl���C�XzSڸV�Afs&Ni��ǝU՗�L��RRN�:���:b�O�H��oP{wS��������U<��j�#4�xK/��B2�t�W�ʒ'X`ͫ��pf��Q
0hf˶��Ǥw��-/�q���a �&��OX7��6���ɾ��|����4g��p>���-5UT]�=3�{O�7���k�����i�n�ѥ`ll�����+��̻Q�ɀ�iWڥ�Z�G�5�(��]`1��Ȩ�t�}��ӣ7˫�T�-�Be-6��S�p��+��)"2x:�P�k�Ju����ﷵ[`N�R���E��_�������T��\� g��,���C^���&b���;��윮ko���F�<k}��H��Y�4i�Jwzx�9`�Yo�����8p�Szw�=�[��<x}0�X5�H��J�E��� �W�f�k��x��x._�)�Ҫ}'�v7�k0n9�x�ѵ��~���1��.%�`n�qk�����U�6T44�>������b��&��*Q+Т�X4�`=b�w�����T1]|�z��Ɂ'����~'8d�ݤl��a�F�\CT��$W��K]Ia�M���R�ϳ�9�^>]���4�a3:T(z�����<̪`
���v˶�a"7/�]:���b�3����[�����\��U��r��7-8g{.����p��ٽ`���/��U�1��0K�n �@�c3 `��ŏAA싟z��45���Lp�ix����Kv��b��l��%����C��:w��}�C���,SV��T��������ƱE��_Ձu<5�S8�/L*��RV喘�t�\���Zc�tӓ����'�M���G��C�"���<R�=��ha�Ѯʹ���K:�����⒒n�ٽ�Q��RH���~�L����wx����!-��o�֜�����qK���ˇ� �Ɔ�C�~�HTn޴��.��g�mLsQY�@}EjRKuU��� ûS�ׇM�H��g���;�I���#Mg���\U?��Ouז�K����D�!SZ��(��t�M�?�B�9xJK����fdd���n�}1����f��f�Z�4���|lаUVFf�{2��qN�}�m��@���.�Ϯ��$�>E�󦴘�}"wϰU��0\I1���F��-G��"�k,��cj�=�^p�I��7���_�'@�����2���I)<��� kZ(�n�<Ң�����F�����>��#���_7K���!� l�����Za�.�lC��5_���x���z�&d�>�y�c�������������v�5f�%[ -�9��a���_�.��N��7���>����kǵޮ�8}e�Ys���rM$GkK58l\xRi:���ɚ�̖6���V�cx�Q�m��7����P%X;��-H�됱7n����`�6Zf�\�!��C|�������?�g�*[nͣ���!�[?�����)�Y^9�T&��6���Be=L��s���YG&6�<-j�FydM��dVj�U�\�"'�4��A ��T����;�
��)5T/~���A�r$�1�2 ��bz�ؽ��t�E�S�2��~>>>'�aj&�[-[ܭ	�]����3@R�����?��kN�]l����.`N�A�������J������I.���Sè!�y��Q�<ב� 󻩡Y�%����I��Y�(�1�6U����f�p��-tC�W$��\2.�(���)��o�&., .ϿϝG���8~3����ni�ؘVg"o������i�3���Q�GK�EC����2�Jj��v
��h��ܬ>xJ7U��aV��<�"��s=��I�r�����|[�6�ܢP���?,(|�}�"9�G$�%�h�����v4`:�w|��&s����󷮆�D6Hayo�������V?EnSH;\�y�zǿ!-�!�qb�y��W��=�k9\HtԒ�
FZ��x.�^�-t�yX�u��3�Byώ��G�c��l}϶�F��l}	 �s���wX�-^�
ZvoB'=u�P�Kn�#J�4U6�^=��$M��%ci���,���?Ev���l��Tϣ��"�E�����|fF����/ŹV"o�����|��Z6qF-����t�I|�`�z?]'�yN{.ęr:�}]����Z^~x�u��������H�I��eѠyvRV=��פ��	�ϭ��!���$�
�?@�[:v�t͙:*���R*PK�C�U�=i������*�'�'$�`�{�/�<%D�]+,TK�qy8�K2e L!��j��>��7�ଡ଼��a���]��YӺ�+�D���i���|Mڝpd��t��>��C��� 9s��kU��g�,,r���x�;
��p�����h�AB3���r��,�U�"+L�Ψ���j�SJ�o���-���{H(Z��W��.�G!�!󙾓#�Fo�7�����&j��I��B��[��ʲN*zg���Ը�J�$��[����ڨWYj���EH�Ѓ�c/��cc�՘s|���X�R��@*�$l��0���.:88��G:�1�z6X�g���'ݾ�e��T�����}�� �`�w.����(y��l�Inl4��;7���������� g'waϻ�j���W�A3�jRgցFB�i&=���	�.�|è&\W�O�6`�&���K.Z�{ʦ�z ��yF-a�`���	��t�Ul�L=����pr�&}��+1�e|߃��CT���]q|��3<}���(s�6ѱo&��C˧�C��["�4;�K��M�����*���$�����U=G���Yɛ���Ri)� D?=!S�(x��eUy�y�1���J��❼�U��ש�:>�p�l(y��p��-
ۆ������ t���JIL�G���D�0�0�\�+W����>�RRR��IZ��A�篊���	mW1*�cO�1鸧p2?��U�'��������͘�U����F��t �!6�8eI�:y��F�����b�m��HD��x����C.��b����f�4�o({���>�yy��b��5��_���H�jOO��n�X�
wn��q,٨|�BA9J�nX�NMV4[�0��^��YK�+d��������²~\7sk͔�P=�Ʃ�y	�����rK��� ���-~y�� �D�[b���q߸���w:��-h$��(�_ٗp�.�J�'d�1yx$w8&Y��Z�V�����%*�[K�O	�.sL��m�N�7��	zض��j����%�"�v4���R����9�6�y�|O�i�ZƆ��I�w�,Z��q�g(�����]���ӓ�4~Aߗao
�Ub����{჌o�n.������_Нx������{6��~?!�,��ս������M����|"?tG�"�nxj�٫�Q-���B8|\V}̏:��M��[�&u[�;��@���<`y>��� Ւ^n^C� W�ɻ.���UuM��F�������b����p��&��H��r���O
����j��s�Cd��g�D��bv�W{7��n+��B�J�8�RH�5 �$�qѧ�U���7�*��O�ϔ[:1�.�7�s�{��ջ�i�3��GW��{s�mp��I#�#���ж��J?�P��������)�I��4*���v�w�[a���{����:]�k8:�~��C��~�V
������sg� Ry饩"%�h(�N��]�Bݱ|�S��S+̨�b��ѥ'��R}�GO'l�GHl�����X	_�l3�O�VZ���?#�6ڌ�<��]�$Ƽ���x�4��Ң�lL[ď�	3F���T�j� ���Z>%Ѽ"��I���KY֍i�(s�a� �����\���]�Õ?l���;Y�����5M���zQ�5w^�p�4]7Q�s���N��~wӽ�jA��@�LC+;��M��C�p�w<3#�8��������V�K'I#���Z����M��uU�������iy�g�a��s�sM��c�h&��R "e]W���!��I:���|?A���/eee�deU+ݗ3cw6��q���EV�D%�~��:�4l���q�ڇ"�-6Ѡ����>D��VM"Tz�!GT��p���`ߣ�����D���,�j�@2�h�`���b��"U;� r����(w绾����Y�N�����r�x'�/6f�/�Z+G���`��W�`aJ�0�tx\�Y!C
�`&�;�R��a��� q����3a��c�����>�*j?���������Kڝ#��XVg�l�3���HU���{�|?�Bggg�I�|���w�}uE����bnkn�O�b=�E�OO~ñO�.y��b�8���Vq�����1u��kb�zo[v�|�Q��c��̄�`���&��δjD���,�659�G���9�zmN%��ܬ�@�;ȄQ\��蹌k<z�� _�Ko���p�G{����|@�sj#����З�;�GټW��&�t�D��9�懝"�S��r�Ϻ�(G�}d�j���/s����.K�\Td��v,��:�r�aP�duNe��2��[G^:}t�Ta�pA��I"]Q�@w��Je�R�V�3�e+7*�O��ټ��9��,|���|s�陼d�>�b�Z�������q����u�i�x��W]S�|v��H���q���J����<~k<�<;���z�(��Ze�SI�k{�&)޲��A�&�m�p�F�.0`�W=�C�Xo���~8���hk���E��9��a��v8`��ߺ�4��d���{^�W�(3���[(��O�hǔ�-衘�~��Wf�dY�R�w��L�$H9[Y*�'=��l�:r�)Ҿ{����y��Rhӭ�%vo�y��|���^�$�Χ�1Ĵ�!(���e��8�a�0]�O�X��nu/���Vz{^�i��z�o}~G����,�r�:�d�0����f�ĳ�eTo�F��^��i�t��~C	@\UD��{�
�an�y���{}u�S��BT��H~1���_�|��M���8�%b�mV����;-^ʸ��?.�X[�a�V`�P�����x�ٗ��e����Q��-w��J��	:����RM���|���|m��#��D�o{�`P;q�E�sܟ?5��%����M=�B=�q0
7�.��|�:T�T���{��/{��.���D^y���(�ı��l����.08�?���p͍�%׶��ϒ�Q���3h�P�U�$R���?e(�g�5��gY,2u�nm�c2�Q���ו�n��n�2S�:
_�	�4�{C��`w��S�;L�;�j�;���q�pP�8�\!�a�K�	���f0�}ɑ����D����,x�O�i�Ɵ�%A��KҒ�}�'S�˿���+�z�+�r�E�6�`�+4yӇ�T�(-��*�t,�Y�!�Z+C��;ql��5i</,I�������v..��̿�z�i�'p[\���H.���0=u/�:����mc��t��P���YV_H�������Q�L3�����^3��&|��"�]0��y[����;}��=�ޢ�ϙ�X$mt�bge�j�mg"1Rʎ�c�7�y/���� +�}ߣl�>��Y�mD�R� u�|aH���\P����_��wj��l�#�U���!'�L�n�*{������dw{-pH=�Ds8?�1L�>��-O\ϧTe�����ӅCƣAm0_��_Cjs�!���p"Y[u�Ov������~����Z�`p�����[�'A-ˡX+���pJc-���݃mO�[��y�U�Uډ"_�x��	�_���lƵb6�� �+�P�6�b�d�^/=��.R�j��ʆ��b���o2-O�4�
nnڣ���E����9����-�A����W�O!퇓2	��hs�´Yo]7Fagŋ��Ө	���z>m�-�)U�����;���d�qE\���F@��������j<�� ���g�I9Ė���qG:cg_B�Ƴ0�ug�j3Dk��!xPiEM����\��޳��B��566���\"�U��w°l�[N�QC1�mo��?7�������>�vv2����u=�D��W�5��$"�bYņu�F��R��T�Ġ՚������憿j�K�~=Ai�V^zړ�^X�ߦ�: B�E]�^����A�%��W �����r��=�D��CoF�+�� Дe��P��@\I�Z(8Xu�Q��'.ʆ�P��i�|M��򰘐{�����x�n擣�����6�=�H9���T�JE�}�[�_���>�:��{�R�������H��`j�=*����64���5ۖ����-��G��˞엛ĨX���|�xR�-+R����yU�+N�{ݤXk_�k��4�Tް��׺���D#ec��d��e�O�	08ݫ�ì��K��X��O+��Yoj�<_ �XK���\�h@���b�炑 Ğ�j���,�@���[�u�8W���o���m]ͳ9���0��+C)7���)�O2Y����{e)���TE�v����4��\IPa�5�5��SW|�W��%� ��uᾅz�<±��N-M���U�fc���..	k��ю��F#:�u����"`�츾Ikx��?��(�M��R�,N�����ӫ�G�`!c��GMƠ�n�u�K��O�/w&�M0����^~�b�iq��UaWQ��\O��m��C	��q}���C>�!?/���$�_V= �i�,�-��~)�ьqF�foYε����$���'��ޑiM�4����Db2�D�����i��pZ+#>pQ!����d����H�M���/��v�^����_��k`H���=�?�Z�o��!c�)�|��O=��ޕt�������M�N���n6�+�����z��Z�d?�Ke���2]�?��"�N(�%���Ӟ�Nw��n],�T���� ���s��]τ5�5L��OuT�w���S�cT�fW�V�@���=���_�5p����
���ë�g�p�x.�)Px龏���nvQ�!�ĉM���Jp���@������eU�S�J�,�  *&y0g��E��q�.���E)����Ѡ'��F[�5SB!Vw�8N�W�)�U��OBa�߁�wr�����:S�����a2B�ge�yT�^�$�}�SH��cT�~+>�s�p�$�um����RZT1a����i�^����}����o{Gr�����'w�^ȃ���hR��%Jh�#�+I��s^�6~Yp���)_����if��I�Vܰ�9��*6�ѭ���z��Ƌ�)H�}/?d��o�̯Q�(Ö����1ߞ���� �[��o�/��u7����#.?�l����B�RP�:
�}����L�6��e�0��~���lwJ���|K;)���| �;Ů�����cGJCr��=FN�������Ө�Sx�,YchNqfZ�n:Mj��X�g��hA��%�}i���d��)K7�î�%��V��h��.K���	.S�I��J�Z9몎��҈۝>�[fw�ŨhOgX�{�xo�vu���SP^\�h���
'	�ٰ�搽w����1Ȕ���r�2tn��[�;���t��2f��gSP�6�߀���.ܲ�-
]��^/���6i�ٻ�]膇r�(_/\�qX����7�4d3���><ġ��!�.�E��k��T�Y�f���ϊ�d"&1�O�/�/z����G��-Hٯ����_G`�Ft�h�� ڡ��3�G�b�Ͼ��wPY���Kͦ������ԘO��+�}��?v�m�0�t$�F�?�5�K}G��F�S��R��[�e�����C �� Wv?5��~>��6ތ���zFr!�,�&�^�E�Ql�>��*u�̋OC+�,_���Bhf[�̘�sÀ���x+�{����(mxe(�<2�&9!ꝎPB��_:������^5j|����7����N��'��N� #�J�k}�Cw��l~��Mf}؛ѵ�������e5{�h�����!�r��K8��۪pVY�%��qK���%���9��a=�.묋�! \����YGE�vPPP���D$��Vb�D��D�z��%�s�i��A�s������u���8g�k�绯�����#���n:*�Jv븖�k�ˉ ��%z��D~|`���#X薰d�a<���u���"��+�uR���iW��j�xI��e��}X~@�!Ni������-�nl�x�l��^�߷AZ���o1�P��x�D]&��� 8�' Y�����yM,'�1��ٱ�����9Q�Y%�KE ��RBi�����ysb a�UV����)�����0�i�E��ݙ�cO�"Q�m�S��H��
��0sy��5?U������Q����ENU��t�aѕԉ��7YO�ML�b��|Y�~�d6YI0C�Wb�8����)ϘL��o|@<Y)�Cj��rA��ŸF��ft`	��֮3n���FMЉ���Ox���.�ӷ*����h����N��2����1HC�]�?��FTs_,v�o�*��������KO[�' ��xtk��h�1��3굸��&�
�e�.;x�����n-:H����
����Z��I1f�F4k7������'B��V��.k�����;=F�i��<ΣD2EE�Ba�E5̃����봢����譫󞌹(1!stҡO�!`���v7��~����]�nu���v�������m�J������=���F��:帱�(@
��ύ q�u��m~,��$OH�Ѐ����6����5?��}R�f8!���#bn� ^�J'�̱͜� i%��.�ۭ?g�5ޘ�6��*K�W�G���d��-ǉP/N��Q��z��#w����5QNF�n@i�4>��ǡ�!����6�w���[h0��l�]��{>Z�D[���v�7�:11QC]����E1a@̜�6�T�����s�ݿ�䥕����?D���L8ӈ�����+�Ƚ��+ݟ��)FT��jMY�ר�q�6�%������ݨ�������PBj :J\�<A��b�o q'i�#9� F���+>+^��� k�����8d�uᮯ��`N��e{�Ûߓ�1���Ľx�千:��eAOͅ��X�[ ���[�E�? �	>"�T�$+y�=	�q�t`7�;6�ݭT�{�Oh���4�V>�f`����v%b�~��!�`���	[R�m���4��H��]�Nek�"�s`�Y���Ǣ`��38P�d��޳*���c/�=*5N��.{7�?!���y�d��4�.���V���ͼ
M��'^�{A�wh/\�"(��s��
$�QIe�L��Sp"��l��x�Θtr$mp+��p9[����.Z�j�U�BӼ�gx�y8�h��I[�5~,����u��(�oal���}G����|oYȋ�&�����h(S�83�T��0�O���Dϟr���y�x�S:y�5��Fu"��]�!����ޅ봗���)�*!{�.ߕ�'y���q]w�?A�	!t:в~ہ�gR�嬉�R��4����3���t�$��[��(כ��!*��v�h(I��B(��5E0�M���}��z��R?��}%4��bHR��/���r�����/Η��5�?.Ϭa�6�,! �Ǡf�v��i"��f(k�L[�4%d��K��ci+H̵ֳ��ܹ�t��#�~q�
7���3w��-iI�)~���qo�2'ׁ^��_d�6Wgd�9?h��y ��7O�3Y,I���)�	u`Q=��ɀ9�z�۫P��Yv�q�&/�@�|���~��孰s�(Mc%%�M��Mr�f�G���'��B��UߞA?��	��R������'3�O�='t��]�n����5��@�/?����I�Hڶ;N�+�A͞�`���Z��o�/�v�i�>ү����Q�^_�2����[�2YVP�ʟ��8<y>�J��P��M	�LK�NyŜ�F)����]�-�K�jQ�O,&�`\曉9����C��>�o��y���3;\�)i����XC���s[Z�nk����k3]ӏΠ�/Y
ύt U�|�ps��������B1���H�*�N"|����$�͆����}&[�J�h�Xat��$e[��	 �F,^zx]�KQ��N���p�&09<@���ŏv_�����=�-�tEl�t_���3^�`�e˕���T9&<��/��Ht����gt��d���p��C�{sP�B��'\�?۝q�s�6h��+�`o�����"��l"RY��-	�> ���.-ɪ(���e�a�$�.���x|�8[���a����&wQ��u�l_�h�H9\?�M��wǔ��F�?��BI[4||j�W��f�|mcMtN!��� ������Q<�~C�W_�S���ȿ�\��P���������~�{[Y�Y+;�����z`%u�ǁ�(]
y94�_L��4���!J������dt��%��;ٓ��'˘���4?f�Z�;P�&����/���H,mI����i��h�j��<sK �,�$�Njj;KPXk�K��Is�nxY*��y8A�o�w�`�
������T�v����(�{(���[.*���_����B���[C��LV+�"�F�ou�.�X֜�~ܠ0����0̬��%OT��.r��D��j;�g��3�v�i�I#r�˖�`��0�':��/I)% F`_dԟ�j6-����5��Wۘ�芌��IN����դ�p+]б=�#U׮Qwx�Ba���rQ�U�w��������~�I��֐�1��Sk.�����wf5~��)�.�R�~+{|���]�'i���i��;[��{~�`!�h)��&��愔j�,�������썱O
%���rW�v0�i�W>����Eׇ͞au�نn�w�S] )ʾ&\��N�@ư�I�܊��=`4Z�wN�N뤁����6�ʢ]�aO�^��4��s �f��\_	��T�<:@uh�z���2��iR}vJ�g_ܽn�:�\�y���A�(����EC��cj&j�zP��[,o���o�Ə�;B�y���`��zH�,�"�����C!��r�r^B�̷*�lQ{Sr�[],O� �fͫ�Wj��'�Ee���y#�����q�3��x�Q��\��R�H��gȗ���}!�{GID`7��i�d�5Z�[��{;R	=�x��&�d���*�V�����.�?\X����{�XY}Ze�]zoo)��V�v�/�n\��#�9��}��Sh�&�MDD�o�}���6Pbv�����藼�"Ym��g��7	�a/�!���U���1*{g���&�e�^9��_�����c��>���{?��#࿀$��ȱ�V��Ϸ�
e�5���n�n<���c�^"D����`yB�!W���~��,�')z�X����}J#C�?�O�]��FoFO6�S>|,C��<�@fT��t�sû����U��H�P��wʄ��52�H7���:���'TT\J:Ź:�[Y��X|�Vx��}����-��͎zOW��`I���C�\��vk}	�bl��NХ&��Z�`�U}�ex����K%o"̔(�G��3h�5_��(.���*'�ؙ��m��yis��U�Nz��_����}���"JkM�=�>{�]H;B�\ܴ_u�zg�r�+���angV��P�p�y��aቜS��K3Ϲ��F ��Z4�p��&�J�eϓ�������7�grXڀ�6�"���Z�.��\ �	,����(���	${f��'�Ϝ��@�19p��_�"�y}�E�u5U-��?���1��8�����J��J�Wy}�ڑؔ�%o�-a�-z���.�F߃���*���:ĝ�u��p��"�25W�PDL(�ԩ�m���8�vO�����$)%�@+Z��j���\���jTsz��ڧN�K��O,�����~g�w�^~��䕕i�В�c�\&�@�u^����E��7��
�X�s���(Et_OU�v���N��ގ7QÝ-��]T	�F<y�4 f۠����Ф��l��kZ��R^��U�0B0�n�ɖ��̀��&mةp�������^
����,�5�+�3:Dc\A�e�4��SX�ڝ�Z*��bhp��͗&���	8XNV���N��ž}��Α�-F�TF�Iξ1ɧ��W5�<�`;#E��	��1���}��3b�1�����Y��kRn(N8���fh	�G:� �u�K
��3�hi�Zg�c��ɜ<��~��a�!��ys�i{�������9������-�õ���jE� �����?B��Y8ۆ()3��G*"<���rA���%���3�hl¹����D:��v�\�ƒS�1�G�2��};���GeeN]���x5�MeX1���NC22
��Vh��?	��S��2��m���c�X�аm�Q��3�4K~(;TN(M=;JNS(t��(n"r�K-͹;OC�Ծ�X��߿���C�dQ7F���� ��W\�H�����{��7�#�x�b�+�Tz;]M�kO�b.���A?�1_l�U[ p6���m��hѷ�0��R@RjLa^�I)��Bp�ۿ����y���a�#�l�}�:9olP���˕��IIn�2�r���;�oKo޴���y�y��j�r�2D�� ��竀�TTt�8�L3�c���C��|�|V󖉱P�:<L��	6B��̀��ǘ/L�~bߢZ�z�p��|j�k��8���64�acc�|����	� �TҶ�vR�}Ĝ�"�q�x��~�h��Z/�;���Lv�z���㹢�J��r�J����y�)��y=$�q�� -�S�I��N�+�m!���J��[�d�+�a�b,�1V�-�.�ȩ>���<���d��E��I~��˫�+��֥�P�,���e�
R����D.��2�\"����L����:@y-�$��߯؝i'#�5m�U �M�͹τN�-�-�h��A��>�~�� �*�K��;=,vn��~ �կ���|-��|/�T���z����x��q�`�څ���Lc������t
�Ϡ�&���Y�p��÷*ę��"�\_�<�c#Vn��*��T!k��2�<����RϳC�2���v�5���s�o***���L�;c�̣���؎��jOSOVݸC��~������͢��;o�%��|V�"�d訶�YH�H��P,ЯjO��K��+�<����V�k��C#�F+��n�sJ�9��Q����/Z��6��h����y
�k��'�%�����
��`��H�1q/�|�Ω��U�B4��3\W:1����|�|������՘��B�Hk5�8f�2��Ff~ajJ���F�6�ފRF�v�{+��j�wIO_�$�g�S�Q�Ƈ.���Q<G�d�Ǥ܍��:Sm�_�!ެI)������_T%iX����-�a�3�$=���" ���v��M�g��_�}[�)��\C��"O�q5����ގ�	��Z��S$0Y��|���I�z�tl�P�Vv�
^��v�Eu�x�د�e��"���p��&c�=�pIl����j�q��:)9�H���|�������\�̈����+7�X��g���f��J�<7�n]Z�ׁ�9��*�w��Z��O}V2��s���k�4����DMY��D��ꆷ$| JA�ɪ�OE�5ԿOO��|�j$u��p#������H�}�(�%���[�
�k�W5
�c%�h�aC��c֨�.�A�Ddِl�e��بb�i��M͘���$�7(S��*&�u5�3���;�FCH�9�j����v�tg%z���c�*|@<9`�����V�lcl8���^�K�)�o(g@,;�n��U�
{�I����*�>Ӂ��Y�Ǵ��(*��m0򹑣g�<��� ��Չy��	y��o�Ab�T��dr�cˈ�<G�H@艐�Z�(���O�6,�D�"뱽t�Ų1�(:��m�p�*C�8n>sn-�`z���v���#D0 �)B�FL=�[ (Շ�&��������i�v��N�n0�����qS����k�,X��e|����+�˟<�ٶ�sN�qV���ꪻ��	{����QɄn�4��t�����<\:��`hx��͔�d��A�R6wT�E�p��7wL��귄
�}RƅK����9��q�{�K����$A$�A�^>=ki�P�{�q� ��uB���' �ڒ/F0�S񕖶n��r)E<�s����/u�f�\
|��QY���b��(_�,�ڨ'�!��#3ڊ�bYbt	��@�h�潥��vn�� �LL�@ƫ����|tOo����XE�3�L��0�O�-j���2%%D8��v����'ҁ��beJq?�F�P(�%�$ۂ�a���[��wk�Q�~�s ������E��־���A=QoW���˄?��K�����T-p�$K(%D����679Đ܋���O��{�� J�N��*QD�Z��e���E���qW��x�3-it�x`�~��Sd�J�ǜ^�0�c�LW=��E�����|�W�N�#�h�S�́;��yi%�Y����� �YH� ]�!���/K?Qz�2 �㄁Tm㛋�G�Z�s��;�!o�b�F]t���l��{��߄t*��ō�Ú���C#�]p�n_U!�J��]��K�_�s�8��:��|b><��?DR����M��Ec,��B��0�IT!�V���Dķ��Ѷ��,?q&������=���K=����V����O��Ԑ!Œ�=\BGύ��e�C��W8Y�X��T �T�
$ҖDi��塣�j{�NU�<'Yˬ:�f{��&��.����c��B�XGIo��/d�wk�2sP��P�pD3�����s"Q��1�Ξ��a�b����ghk�n��ǟn/���ݪ���-"5l�0Y9WO����?�T��Ud�����2w���ȝ�����տ.�%�޼����VB .�PS����Ѭ��+�py�U)�G�����nw%^��{�c`:�\{>~��X�B���c̯`�>�M+ � �C{��4IK��J�q �t^�xx"%Չ�6 �� ��+ �˭̺s��#)��s#^�w|�!+�hj���?���]鎿W_bx��y������ө�Ҏ��P\��%(f'jP��=O���L%x4�o�O��<���yO�ki��D�����D	O3��no���� �
��%����R��eP �#�{p����E�NJMz�]7ϟ�ȃ��ؼ�N�e��+�:�4Œ��Is+U��̞᷆'�ҖM,��;��	6P�B�����w��< X���L�����3z�Z`��*
����o�3|A;���*7��K���y������ԛ+� ����7+q����{�F.£�Z���� �;�R�H�(ݍ-�|�G�7y	�lxt$҉���� i Y���ѵ����[>	�M��ݛ�)KKS��!YY?1��U"FP��G�=�}1<K�`>}.�C VxUUU�$&������.�Cr��P�ť%���c��1�.)Y��&+��$�?!4B��a��>�"r�Ya��!�[��[�&Ե�����B���GB�=��9_�>��W��U���ۭ�q�M�P�L�v[l�^�p���HUYY���l��#3c����s�=T��� �9���-#��U�J�w��0s,�w{Y�FP)�.�M1W��2�Ey����� �b�.�X^�8���_��7(����jj_���32ީ��g\E5�����R$<1���żB[ww�#{Y�Nڼ�\�J,��ç|���������|&�'X�d|�wM���
��k���U'pK�����_t�c�>F��M<[��#��M�r�߬' ��M���~�)//��2lL;W-��񙙙-.,t�#��8��HC��6���M�74[4�L	�XVd������[B]�W���1�G�!�\.x ��8����Y!��?�gr�}��%n/���?�b�K���L�6ft`x8gc����#r�0T/N���,�����0�E)#\�G���7J��ĸ���c����;��o�L��x~�;��]fϚ��� y�f�+���hzWB�)�+��D{��=�{�C[e_U�ߌqp{���Juy�&�\G"�4>H� � s�6��M�,L�Nf'������ܡ���(�CE_R��8�_�3҈GxB7G���5��8$�/O^��w��,��24,(Я�Ō����Jv�څ�YvЊݹsG�e��j���2'�k�mz;'^�׽"��<;��F�9<�� �@���(�ă�wk�TZ��=R���Y��i�'�Hj@\�k��v<���F�Rv=@"�rso�󖔆��B���󛗻�}Y(�r�QU���5[S-�isvk"��a��d���Wz���N�Z���N6��*yƈ>��N�cPf��S��e��Tf
u��υ�X��V�f��p��=C)Y��ڶ`�Z�o߾�{���$�.2;�O\2W&��m�C1$�_��r��n(4�H�N��:6G��I����k J���<�3��z ������Sx��|�|V�B� �i�(�wՔ�N�\wwD�ȋ�#�����Ec����8�0X���;����M��ubc��J8і�"��g���(�����qU X��r1�b�ݼ���/�%�=
wz_����e�����Uθ�B�*��`k6�������M'~N_;�V����F��f�ᅅ��/8ئ����j��ǼN���R�LW�3����_T��:o\|�j�rdN�e�<���g����ڭ%�R �cD�<e�`_���X~`�dI���Tmބ#��	U�v�_D�=W+��N��s|��g��E�οug3ipGݭx�,v�I�^�v�����A||�'��Z*���H���Cn2��Y;RjNKG�n�W�j�,)���Rnkk��!��<��p��&��i^��D�#m��W���h���T�O��D����?|>s%C�ߏ�xC[���x��2餛����Y�;�V�����կe���|&z���{(5xg�|\j�e�U�A�6�".t�������Oo��r��`�nBy��
:7�_��	��@��o�a�ݓ7�.�������8���ge��Be���bFD���\�|~��6�@O`���tCC	O߈�t��o�+	{��
S1�8:�(�����]�n��B�_�Qd�ϲ���֌�-"���*]p"�6IR`aV	^�C�>;��=��:�S ��f<�GG���Y������O�<9�֛�_C��_�B��$�r#.�I!	C��Vb0����I�Jk�v�`������98�IQ���c5�����4�����E%�wc>F�'�}�>�UW����	��,��u�^�t��x��9Ÿ�P\�*!��ˎD+�UV=N�[;(��lǫ\���÷��
'?Ì������"���NV9Һ�\K��n+�@,�r؝��,�����U�eQ����N��(c{�\����c�+�����5c K�+�Yd\g\r���p����RZ���Xw���Ķ�\�)�WQC���t��qZ�M�7t�r�D���J��)�c�,���$����MYU�ߩ['��Zl8-@-�D_�0'}�,���w[�~�w� 7��h�7�p�ͪ9�Ӎ�����~���6�1�	,vI~��e��F�M7�(��������@fKmNS���$F�kk˨�3�0�t?��j���xf��p�J�����&�Z�_�H��� � 6�ݘ�X��=v�c����]��%���?�m��
NS����}��^���'v�T�4�K��I�S�lP���W#8�����gY�x<���>���/�s+�c-G��`'�<>��v3����	~z�n�j���d]�c�ͭ�40�;� �@TR x8�U=�\��Ȟ����������	Е\@٫��@��jb.��܆��^ ɿ�_7��Z��<��5�3���#�a��7>ON���MK�u�&�����=�v���PE��������顇A�b�y���J�	�%,��\6}����g,�q��dgn�}����3f֭���M�q�ۯ�wJ޿�x�j���A�:%h3��d�ʱ;/2�G�a���9a�Ƹp~�\Tt_{�g˺�����w�����d��`-ǥ/^�Bצ�99�=<<~wt�l��Nt�2�3�3'EF�mn�ZXY�[IB������,�I� 
�ߚ�F ���l���+D��Q�P�v�%4�
=X�\�&��E����Zn_�{�:����xj��7� 33x8�1��I!<S���K�����ǻ>Qe������Ģ�����ú:I��~P�w�R��sәOqqKQ�\ŌLPﭝ�<�8�^ T8��	H�˿ ^����ݚ����_{��V���/��ߧ!r�|{;\Po�d�ɯ��� `�Y��YHx7�8�=	l��ޝO-�s�|8�.�8�0�
6������_*���D��q��� 0�Z����n�s�7�Ȕc��HNN&z(>�k��z,ՍqU�O>T��s���^h=Q�sb�a���}�^>����XP$��f_����3�8N3׹��_���A�����?�b@ s���A�M�=wk�4"%vO1va��ٟ������oֶ/��X������u���X���J;��{w}6��t�e���X�Ų@g�P�Jb�z��#CL�r�G����#I�{>�8� �o-ĸ?�i����_!4KX�ʠ�*]���Kd��[y����!�k�(7$�/����d����nX����&��"���c��<4��3��M <�����a��%��b�g}����hq�^9�^rG��,�ql�n��W1��TTy-�}:�?)U>zxͧx�����(ϥ���o��p��R~uQ�FF)����=�{�)|Mf��n�+)--��Tja("uy�7�1�K�	h��:�~��m�c�@����L�^�
�F��ehD��{�M�)��~��ϲ=�q���H�Ш +�WOؗ+�Ͷ�0�o�fi%Ǥ?�9�9�&�yK i(*���<v�Q�a����z�D�F���MZ1��{�(B+�܏����ť �M]T� ��P��粒n���G9�W6ga��k�=��mԡ}Կ�B���.?x�" 1����}��R����*����aG��GR�S�;�U��%k���[��+:E9����Rx������q�M���V�Q �_����ո�o^0��}]����+��Se���4<�'��n��L�H���6�>G2t<��K\�=���K�Tj������DZB9`�L~v$	� ~J�JBB�:�kv��06N���x�H�4\��+h❙�V�z�|o��d-9�~E�OT����7Y��k��������>\��I˜g�π�5K�~���PZ��B�@8����ݧz����lC�U�����rq{ԩ"̢ϕ��9���s���΂��[X��+*��ɕ���S��	m����o�쬬�;u;�ze��+����l��ֳ6;X��W��Bh��\�_�d�)+/���y�Z�XTC(*�l��z-~�o����4�}���{����p~}.],����dݰ9�v౔�W��بk��&n����_��
�VͧT�����t�7���,A/��"c���rG���E����-p����a�A�������j�Q\�����Ǡ���uw6n����I��<��r����J���ԯ�wi.����6����$`�����3�њ���n�'Yj-������^:�g��� ] g>.O�G����];�zӟ��NtH<��;Ԯ@A���D����踸,�ѵ&�Ā������D���v<N �>s��8ލ�孰TZe�n˙�Eb��`�C��� ϔڟ���wnm
��Y���}�,���I�����<8�?�w�u;�}-����c�M7�Zf��	����TT����iT��?�m�xc��9y5�xg*�C[��焏��%�!���棥F�N(����tiS���Ǜ�c���[	��j�W۱B���nF�l�v�:���l��;"U1��<X��@�Qf/�?�.�a�~����@N�4���rk����[�+b���H�[��Tj{��w{�%�Y�ѓ�*z��P.���<�3֞{p
�5��H���SA��1�x¥�'ll=;�\�:;��|�z.Ѯp0SCCG'�[�����L��b�~����؄���-�gFAQ�`kNE�.��.U�w�� ���J"����q�ۇ$��� a���,�ޑP����6��u��xя+W��sssJ�V������t�n޸�N|�Ӯ�xɮFO{Z]�J��GTi�|k��Eɮ�OK���^���t���>վ�rkjާFE]ů���� ��[\��xo�K,� �S�DQ���6:Th,�k2xO:V]-ڑ��\M��4m6^�1R�����fm������1C,jE�~�����?�̾L�SݦN����~��B�T�wy���<7���m��	��
�wp��"�>7�
��b�7�a6=�}B�V�S���5+�Ƈ{��h��G�ѭ]@��[v$f�~Mt/I�� ��i���y��ZU������cK�'�{&���r����W;U�Y�o�4�
�L�,�aD�2�^�~T�k��ǃ��!*�%ZlC%�/�Q��X=ߜD�˙�� r���+B��\�ki��'&%�������C�f����'o��]�,�� g;Rf� ��+G��`�Z���WW�t_��R;�sJf%�۠��,+��n4�P�(�T�7�P��Ӓ�)�:Q�Z%Z>k�7QY)2�'������>Q�|��а�	&��WM7J�P:�/�����>e�_��������W惃8�U>_Bj��'	xK�j*ٖ8}7Q���|���g��n>vvń�����]��YRܿ^h���	��0@����^�g�/]��.s}E=i"{�
8�[�|90vw8Qp�I��e�J��"�61�D����+1�������"�nB�}��~���J�/��L��1~�"��V��s��?�!>��$��%�A�l>w6|������3�0���ʽ׭�uw�'�Zf�,�������oI�e�����nN��KnvvC����h�{c�Y��89{/O�M "�{�|p�6z�5Wp�F�k�x�>�H���qo�E�~x�1>�?^�������]I��6����g��^G�B�F������*�p�҃�ٿJiUDf��+ (�t�r����Z����ʞ�AJv��l�vP���Ez����Z����C)$��+kO�R|KC	h����8B4t���U�=:,_�	�ѳb��(�1��;�WP�3���D���L\<Y��V�%+)\�@���Bb��Ӹ8
2� Ov})LiΞ��󆂼��[�$'�y��?�O���r����(��eo�;��7l[(�� ���]<5J�����C.I�^�<����/\T877Q� �
�G�����juR�k��p���:	��"�[�r�b���^�T���oQV������յS�s�Y���Л���QVn�wi\j�~��w$ku����S`���]�o�j�[��B�뛳*���Z܎%�4/�w[���e��j.�&��[�� �X=��K\n/+��o�i��ɋ?1*Ԧ_���42V���yT�Ld��<�&���5�(,���O�V�1�W���_�퐹�ᱝ�ׂ�����j���׫�S��Y� Ps���;�t���7��Q����i&v���)��'v��+|Tl��av��9f��(���
&T�2@�w�l�Glc۹�?3z���e�OX`Bn���2�� ٦\fen�9���8xqbDd����7�
�pF����5��G�������J��h��ڊ���-��f&$��V��~9��o������[��@���^T�s_�B��OG���!鲔~�c9-�K|CI$y��ED���"����6�Np=��&����g��J�w7�~[T&���yzcb�{����7� z/��� �CpyM���/́e��i�uoY�*��<��� �h����9���r?i;�G��U����%��FF�厣c�2 λ�~;�J��⻃������_cص����X/_XЮߋIq�����
�%|����}�8CHBy��8����w6�}��y��0س��##z���+5�D�2_ x9��9t.	�x��|���7�KU:�+Ze�r�/���>�� ����Ϣ]�3EN � ���}=�n��W��+���[�����]TH���p�j�d���-��C�CΕ����o���Z����W�+Ϙ#�z����(v8ݚ�V�O��T����f�ߟ����IN�D$�{� ��U�`-\f
Lt���or��M9��r��ݶ��)����())������o����x�.�Kq�Oy M�'�����p~��k����>��B�R6��l�o��hM��+C�d��,޵�k��AK��'�uE��֩������Du9�A����1s���?1 \�z��O���'��F@
c��+�bصw*�� ̈�0�w$��]�NE��a�,���,�`��*�]��kbb�Y܃�} ���O��&����2�At���C�{C�XK��[�""���jev�s[��h~2��R��M��:hk���o�*���4/o(��a�(�b�
]�1Jy�6��9�L.���Ҡ:�q��{���>l�e�v��a�~�U���(<�Kr�rq)�p��f�mk#�� ��<�@��t����8w��ݫ=�ܵ�+Qs��xF����GK�gɢ�`�_�?o��z7g)b(<�*�����j���ݙ�.�<�^��?�LiL�c	���m���	�N�鴃pR	t�:��&��}5e:l�\��!�3��<����x�i'-��f��4Hů�]�@�lw#�Yr����z���o?���۳�O��w�?�>�����-GF����ཱུ�ƭ�w�ԏy�`�ˮ5��E:�T@z�G��N$l��B�W�~3pr�pB�E��Bd��}�e��ш�imYNm���ۧ�PZ�(����8��t�vB�u��\���:��v,t�m����v�8���w��~l���%��.ME�D�P_&�d�>�~�+�t�ǌ �y7�Z��x;f�wU�H*�"�7�uo��v�$�����k�̕��I;���z`����V�Ф��\�YK�b�;U��l�!+K7���ꄦIj);'T�KGP�Pt�/�ǀK�Z��� �W�C�m�zllUu�h���&�eė�	���zF���� �p1�����`0T�O��(F�$��z�*��ȔL��P&�K/ᑬz��sV��]��.
������c>i�/����+Wz�j¨<�v��4�"E�6
L��>d_p��+�:�F�.St}�  vq���^��D702�k~��Y�F2���a]�ԡ7ᛇ�t|uC�����^��}� 3J-�A�;R����]p��>��
�ut�ϒ�4���^Cu�|Np����?ä��XX���R.��E��v��Q:�
r��T'u{i&��p�~v/0on�Q_c�hҫ�ZY��MMM�?��qidt�`n�#��U��=x,�Fm����x� N�}7����Y��>xT����h�]		��u~ !D���R��[V�:ո�S�_)λ�=��~�QϮ/��Ƿ�@�۠]�):Uv�*
����a���ȮaqK쥕0![3�C��AM\Y]S�����Ƿgn�ĿD�8
U��Lm%�{���io������8�O��OEC�	�D �4�j̤��`�^��BϷyq�pf�x���C���W��9�����HJ\���O櫘�z)# �����D���P�R��;�d�mn��Sc��m"ģ��}�;�ϵ �t` ��x�����c�*�(z�C�8Wm��(5H�R�$x(��<��{�َ�zTPժ�ր�[�,�}1���,�޼�Л��!20.	��"{1zLe���w-�2����l��G\�_ùY��̤ٜ��IU�,B�����reŃY����$�*��P��d�w�^������m
����擡lRR�`��?�&�>���?�~\�e�$C��r��έ�{������^��ʲqrj��G����K�k�e�O���Y��O�R�!�/�<�o�n�#�7.6�nq(��!�wU�
|��H�a�=!v����R�"��w �i�,,�OՊ����|���E�G����=�B��?�O
;h,vpi\�]���T��MK{��z5����o�A�~SSS�Y�^�.�$8
�g�佧�BE\2��^d�,�� ���f���ԝ�rǏ�H
�1T��Wy)/��0LW|0��\�ͬ*�� j�jInvv?���`5���o�;q�q��t��;�"�=��+�`8K��g\.���Y4y,��e��(�G�C�O��� �����Hz�����)��[�;�[>�t�]~.�ο�I^ ��|�X�A"�/޷�`oIf�P����c>}b}��Y���`�s'�B��0?�<��Ap��r�|�C��7_ә�ժբ��B}I^�{U�[����>���)�`G�Շ���r|�qK�Χ��]��*��0�� |�Ɣ}��3IR���䊎�B�K��0�S~am���ka{�I[�]a�	��~2��/`�~�d�(�o ������������e����Vn�P��V�w*dֵ�"��K����V��k2J�3�.!��I�;�]��p��yfa#8�t!�>���/�}Gu��(�A!yu����K]��N�t�c�`�>�í<�Ӝ]�����6gB5���(u�>�z�k,�& M_~�o�����/;V�'c�d�=�8Cr�j�#
��?�88!���5300���G�&��'�8�=\j�����T�ٱ�k��Ơ�1�og���:���B(�� ���p�  �{���xT���ճ�Sn�,������;F��'�J�rD�Z·e%9���Om�1U��������x�h�����[�ɽ�������L夷y�qX�
��~��8V��Կ�u��4��K�ܯ_e���uK��K�MyO�fceU�������y$���f�����ߤ|��^���*��WF��\C�ժ�wS�Ή�[���n:-U�uZy1�}����R�WC71gW�*Q;�[�7�#�[P��a>r��w�N����1��7~�����~� �o<��4!�V4�-��b�g$��y�KD㕉'Y�Ŏ(Q���~��'倔�4�ְY�Ն�+�L��SR����-���(W�2���YQ�㳾�Z��4Dq���N||~���T�a˚��'Ƥb�?~�� �f;�.�jŰ���U8<��{��@\�]�N8aO\�c��4�T�	$��+�L��p�nYP1���%�ʼoR6(_��2D@.��UU閗�����C���Bc'Nų7E@�Y���鬈���$���'�%�gb�ƶR��z͒v[����=f���Ļ���k�`�#Q'K���w��������hhT��x���n��g�V=k���`�/����ǧ���5 ��b�T����ʸ����AJ,DP,BPiP@@Rj��z�RA:��F�[Z��;�c�{����y^�F�{��{���g�����<��$��͞�����y_��ő�d*.�k�z4�S~7�����7[�=]E�1u��5�ɋ�0�B\MuP	�b�OJ��IJ���tߧ�.���x�eh�hwg�|}L�N�y����^K!����J�%5�b#%%�؀"��fi�k�	7�	� N�wep$_���؉�D(�|:�?�����0`�Q}�2���y,M���4�B�~���Bַq���r?�Y���] �@+oհel���)�Ֆ8cM�����{�<6�7�\Jz���!��rrr��@���&V����[�#X@"���.w�EL����q�D���D�C��D�	t9{�@aD�4X�����%��A��o���z�{6�-s��	S-���#B��t��C�5�j�<}o�8D6�i���`��gх���ܕ�����q�qv�y��/��A��	�4&�����,���gfX澦�����Z�B�����f�����B���5��b��
-[W&1���Z]����Y�����?��r.�\�)� ��4G;��ώ�x`z	I����ݜ�X��Ǌ��~	�[[?�s�Wll,]sm��1�9��Ҁc�>�M��[����yu��^R�[���LO툮ЩetĘw��7��� a�@'���
?��8O�kQ+@��;�u�'_I^�sִ��I� b�+���'qÁ��F�����Z2��Z����zy������[]h�������hnj�X}���G�㊼\�K9�.&��m���y� i��6Tb�"��z5xd���k%{����~	v�SkG�/Ⱦ�̝�>��;L,�;錢)6��.E%f�o%�&.%b��g���(ԃ|����e�@���W$��]��ZB�����_0�yV�
�顃���ʔ��N˳M��\�e�ʇ	��MS�ͬ�E��۬�9��6��#D���Ο���d��ڻ ����uϴx狗7�&Ltur��������GsaO �M�����U�D8d�{�n��9��JpS�C `����\>��6�_n��N�[�[)�uyo�w۩O�r��d���qwA
�x�X��P+�[6��@6(�|�4rTq6r4a�gr�����|��I��B6rj��)�ߣ�~���	�$���z6��38�Exo_1hk�������r��M���ڍ�l�|��X���>"Td9�S2h�A�����@��F��#s��K6#��������	uR�.j{ۜ]f�o����?��P�H��T>7,�I�qNv�-�硡�뫫?��?J�p���S�����,��I!S4�f���o,d�w��{~>A(���˄B�@�)	SUf2��G5���^�~G�|�1������
n0�������yN�s���/�m��e�Y�=�71�Y��t'�����q���>��>TL�o"R���v]%����L�+q���o7���R6>3繌�<�(���������hIT������g�v�!�H�Wr1����E+�obh��I +���!q�\:1��_.P��ޙ�6gg�� ��j��d:+--�4W��#%�)�_3}8�91==h[����M�R��&3ټ_��e���|Z�s���|{���	���t�T�<G���]܈�ׇi/��է�xu=;��2���R.��O��"��Q�Gc	ꛡ!�c��z������TI2;��10$g?��K�U�p��$.,��e�Ӟ�7*3��V�X݅xF��uz�\�te�Ǜ���v����՞?�Z!�{=�����>�lE�l�#<ސU��J5���H�|t	[ff��B�YR%B����(5//���%�X��ó+���J0�uCP�K��/L]Fd���WsP���x~��46�m'�Y�|��/mǪf^6�w*܏N��;kJ%;��|�m�[����G�Gi��Rc���rPK�»No�N}m�9a�zdK	�)'�˜���ؽR��L�m?�m�̝�}~�g�Uh�v[�ic���,�#���Q�������"H���G�q�ݖ(n�W�?$VPWO+�S>A����l�������M�w'D���(d�e��>v6+"��$)�HV�:飗y�A�eW��P}����N1��Q��;ƴ�eS�Vf�k9ee�ttt����yy��q��{nZy��	���$��M����D9��5�HJvg헀H�ͪd��}�����I�k�C;ԉ�φO��36�M�.03��>6��O�9�K���6����.r�1���W�>�oDRu���-��Ó�-5��DAʤ�cw-�)R�H o��)�����J����dqަ	,C��y�\���gl�Ь�m�h�{���������i��IX~���ȷzՋ}�+�z�� �ݘU�B�\���uj��=
b;iǋ����<�c�7o�����B�^W�3	�b��K�
�לl92��|��z�l�L����C磼���G��k+�;�ǻUp�&a���D( lQ���V�q�n��U?�4Uأ&��X	��zf&����ơߥ�Qt\GL�o����*��}i|��%W�&��~)m��2�-	��M�E#�+�>�K,�b��"�cm �:62��*�'�H��He�B�3�]6������!\_�>@��댰uK#5տ0,]�8xѱ�⿽"HZ�!ر|�+�gw����槷zzȄ�DP����t�W�3WF;W��߰�/h[/���&<E������[�0X�p�4(T}tYGI�8����6g��}��|cN?3l35@�F����G�6�H^��Ic*���/pqq���>~3Pd�Gp\�[�@�ҟ�|����xf�bdׇ�b��[e�������	���#=�{������d?w�B�� ?�������0��Ƴ�>��@@�z:xS�����^�Q_����U��Tr�4�R�%@��Ե�?�Vv"}3�i�c)2��X ,m���?��D���z��4ki<�����Z�A��q@5�%O�@~ܐ�X+�y�I\��hͤ0#$g����ٺ������� O�\>s�xdB��*�WPZ����������Z�q�9����ܶ�^O�9�-N�_�F�'��J��L����s�G��F�!;f��J{V&�	��!�<=���S�3��	��"j��V��<�|�}=�GQ��S��5Sn�0������k�*_˨�`����8B�L�2zp�BMH���*��3bn���	N����|#��|\��O��a����P�e�-��.V�0���f�^�>��	$7{h?�����]�b�S8O�B���?9�?�\��
wĀ5���G�
m)BrJP�,u����>x��-�eaQ�r�}}2�Q�%��Ky����k�]��b����+��fM������}I2D�����������o�mh|<�Ȩ��`���`[��ZQ@�G��}%U�ۓF[=��sU$O:���k���z�҅6[����ר���5�]Z�''�&�<|磑ɰ���W(�r������a�>�>y�;�d�#z�� `��2�@~w��=պ�����r[�4���z�����]�fw��=����c�t�(ҭ?a���x[y��ε7���P|�S�n_��ބ�Ax�	l<5�悯�''��;7�K'TA.��ѥ๦bk[���L766n�ƛb��B�L�������<ZL*~|������1��9b��x}u�B�}P���v�q�h�J�Ec��l�`E����'�û&�,�]�uL���fi�O`�����<�ǈ��Cע���� �.��牧0��/L+ NE���;��V�z�c��O��O)��j�.�B�Wd{G�񯜟�KSP(��C�O�3MU\��N��ib��)е?^�����d/����������W$�@>O_)�A�; 1�1d�j��wB�6J8��2�L�Kzτ�x@�:î����h�(�Wo��Z�9o�9^~�2��1�����au^�!�hȜz����O�JS�t����bII�РOoE�H�>�0� ,��W�\�w��	"Wf�d�;����z~�Sw[�M��[Vm�#��ՠ@|�%�>ucY�LBWt_7���Of2��M涄EDTe�u�y{&$_	O,w
�;��U:W����j-�s�U�-ˍ���0Ү�<	V_�<�=������bم������ƒk�y8DtcTZm?yg�TT���T!����6S��|�M��+|��6�ɰv���l�NJh7���S��i�ٳA���cJC���>ldy�Pc+]����$����7���n�`���'3\&M��)q��9D��LI����p_���@�\��m�l�W��$�({���x��p�뭐l�vp6<�/ Z���$ۣ���cvq"�n����v�����D=ku��fc`c��b��O
���@�;сB�B��	?��ePjZg�i��s��9�$�s�0�x��D����Pϥgs��D�=)�khd�F�C�T���l����%���}�k}"����zuSi3l�ꍿ�-���OuS�k=+#}��lo�
nDBWZ�97���&��n���"�W(=�����Q������������˂%f���V�JY��wd8��
x�}=�~܇�1L���y���Bx���畻��x�]�G�G}v�E���<�?�\�I���z8�\'
�}�tp�o�H*�"*U��4�hx�2�~��,4Yw��X�r|]��Xd�]/�7�(��]�FѪ�y���ײ��p*c�V?�+C�	T|9J��m�� l�����~����>�B��i������⥮m��Σ"������ ��[ļ
g��R�+�����ج�
��_�ѭf�K�)kJM�N� �Lci1����k8�������W<�d��⒘�MN,���IcW��F����6���9B%�
�������i�톪m��SH�z6Au�-S����ԛ��\sŀ�c�|�-n�9A��=un�ߘ5�����;5���*�֕����K���;*l��t�8�ֆ7���'�����÷9&:���Ó�ۤ�*����&���01����wKI�1Gvt����x.�0#�=xm�k��)��O� ���7/,<y��|w~bZ��f����+��ť���(��w���.��`�<}�D�@�jbo,�#u��|%�c�K��Ԅ U�oF�?���؂:\�d)�/#�+h�KÈ�7Y~1M��s*�t"3��5��z���^_�(1{hkQ����ك�"]m�G��p-X���l{�Gz_9�⠃*��"D�ѡ�?�o)��.��=vY}Cc�ec��`�'��/���r��2��a�����H:��8�&�#��� Nf	�XU��K�B�4��%���qADF�ozj#��7�sp}&ti?=��%����X�_#j��Cr�,�z����pɓ��̃�i��Vf�bt�o_+�o��0LE�l��6��u嵍T�h[5�W�}Ƽ�EQ�dW~>�̛���+�ZN��	܄����n&\̫��"7w_ʦ�lL,�8�Q�Ǭ$H�Xe��9�������f��푄�ξ��?|e�6�4m�o��]#�v[��ɣW���-�͏�< ���������Ԕ��i[���dś��v�}#������fw~޵s7��!�  �
��q�vS�Tu#�I���W������3C��շ�I��˪K�X�
/h��&�������^�迵P��\:��=��� (I|�j����2�V臌[�?d?��o���ex��K��v��ɼ]|p�=��\?T��5�'%��c�����ʪ��O�AP_9�*������<~X�AM
&�~��c"3�C��#/O��P_�4�_|H��1���t�f�K�?)�� ��۽�(#⟉s��%�@Xˉ����0��WS�������s3��Q��/�N.������G��)�f"<��a�� ɵ*�$�:��J:2�3cKe��e��͋��B$#��SK�N�k�AZox ���{��WEO3$A\}
�VG�(-�(���m�YM�Fz����y���'�:E|o���y����O���W�UY#���xn�V��Τ�RC>�ˡV>{�\��q{lŭr�b����������˧�L�ʒ����]���Y�aTںp�M�+DD�7�UV��_(+�g��w�2m��W 1�z��:��w���`8�R$@6�%ڸýPw�� x/��Z5��A#TY��j�Q�1�g�;xu���M,A��Z������K�j�� _������:*R}S���U@�M��P�
��<OK��tP�M�bQA����W���e'lo-].Y��RY�����[i�sP��޽�D�(_��v!���_����� M�ʗa�����w[_������厞�_!O3�zt$����HݩR��\a�`3���������G�e�������ja��w�?��DI� �l$
�eF�#L��-__b���k����g<�D�x��>j�����mr��Q��y>�����˫�:;KZ:i��O/��$��uz�9~(��eN �V�DRN�'( ��U�oѼ�M���ei�k�&�������osIv9������ǖ�fY�ŀ�11�_��呿`s�Z$[W�ʓ�S?�tW�80hD��$~(F�P��Y�)b�q���7��@m�H��?�Ŧ�����#�P޹��h<��|`�4��`\��k��<Jr{9Z�Jm����ė���o������p�#}mU�D��f��b�Ҧ	d��겤���N�L?b@@J*{
�Q�#��.���-����q��_��&�����,��hL趻�����wqy���.P`x�:�,,S[�4������}��%�!-N.q��s;m�^��ҿwVH]��L`��̇c��5�K����y�2_����|�����y���ƅ���wk�قvkmM��4c��k��P7�H��c�i�KLx�OCv��Z�s-�?>�b؇����['�v�' ;���+��"Y��?�ߏii�u����nv�Aw�I��]��j��D����W���?���`���&��7;��o��91�:�L�,~����M��84p�\;y�-��G�kM9N�{��;x��?�z7���xD��i���s�� ��*��)�O� w��I����Mŷ2�~�O�������i�2��?/?�	++����!v�^��By��
����j�������1��X̉R�	ac˰?�'�Zzbd43�ED���c.����[P�_*?�|�xF0H�kv~�^�`��(�8v�X5#<"�[�f�&j&4�̢�_~�9;^k$is�mx����djJ���D�%j}}]z�ut0��y4��܃Pj�(����5�`�\��N��A�q�3�����{й��|��Fzh�Y�xz����b`�|Í̔��l�T&Mg��;Qi��>����� ���{N��\y�!�NNNm�.�|!l[ABB��o���	�
����vt��9������������uz��O������@e���ܜZ;:��+є��c���W�����9ϓQt����M�u?,�Mut��ee��A��	ק��u�����<PgZ�!��6|=��>(!�/ΌZ�b�����yx*�ڮ���|�� ��1GF5P��E���\����o�{� )�x ���Mߞ籡���b�WB�k�-\���ɜd��5F��W@2Aȣ�9��Z��
�uL+`Amr�7�QP����-�d�Ecfzzvao��3�t����Y&��Z��C��]HC㚭�Ȱ��Ìݵ�z"W�i��9S�ѝ�o�����2�/�q\�����#�}�K��覥��|��_�[�:�U8��"�~ֶL�xjֵ�]���[��1>���6�~��������N�
QL=د�m�o��Y��&7y�`ie� ������6鸓�PU�ϼSc��IOO/�t��?8�X�t��}{�~z�۟G�U�r����B���`�j�kթ2W����`��2�}�Բ���(����J5&���)����u�F�`.nv������>G�zĒq ���8l�����0+�N:Bm��l��&�?tt��p\v��9g`+�D�8�r� ���f���-uU{"�{�du���ƫ5}_�^���3����I�g�����	����z&���s�kक�{i��Y���Q~ĥc���^��]�����c����t\�M��
M9t�I�2wvlyuww���D%�%���P�x�b}ss�w�˷U��9�O���9���OE�`?}Q�D]}�GN�E��H4D	�p�>L$�6U�Z��ųֆ\i�q���=0�@��$��0��$_��r�h�-[b��=f����"����b��.j����r(D4:(���/�i�qu:�c�w/2���x�Aal���-����ǘ�ݘ��K�'/
�.����aL!��<����<6�G`yLi�|����� �«-�ǏEEN�{�$��q�<@���N�Zd
���m��7�K��|�2+�z�����;���Ϟ�k�< � 3�@Ba�6Va��F�W56N��ٴ$�y�Q�4�L#r��M;����b�zmg��|,�fe����)/���jF�[ޞ4�4Ho�g�{�+ qx����܊�}յ�����/���j.Ao��{���ɞ�\`�����|�f�fq�����j�f���������|S�	NAE�����;�@��ϱuD=`;ʣ��<����Ħ @����|�r\����׳!�x:�M1	ɒC坮���x!��S`?�l�j��E�D�D�F"��j��[������.$�<5�Ր�FŸ��{��*���� ���������R�,� o'l����D`{���D��֝;3�ҴE�,�G�ӻ��__n� [b�;
�Ŗ�{��\�F�A�e�൫�m�9�L���Ѷ>�^`��m)���s�1����b���{���	ŋ��n��:�>=Bp(�3�x�mk�y���Ӏ�`ԙ�,�d�Z\���Ą��R8��ۀ�D��z�/MA��h���Q��}�|`�^�ūƞ��^+��yaQ�0��Ⱥ�_TUUUysG�޻T�)B�'�摵5[��/wX��d���h�Ϭ�~4�&��P�磛�9΅�����6T0x|�`�e��D>�cTG����DE}g�R備���dT���K:��u\}���:�l��[	B�3[��h2>�d��F+�cM�v�?ܟt|y�~�|<���i���_p��-�j�vf4r�iN*į>�N�W��6�2LD=22p݆o���\g}{��)��®箝���]�+崃�0b
Z�9�Pq��z���P��>����6R22������/�h�#<�OX���ת*My�ƅj;��<�:ݕd���F\�`������l��(Ee�'�'� =9�	�������\o6|ܴ�]iqܼ�RSV��\�m���i�S��) ���^�ʞ�x�go��ٟ_��;���$ݼ�w(����^=ǗV����\�blBD��(�reO���
+��Ǹ؍$�FX����_^J9-�i����v&W1�2����:+@a�$$�����[�4X>"��:��������N����J�/�<�6�������(P߈M###����~lll(���CB�?��|��]�*��e+�L*����$|�&T?��拌|��Ϲ��AB)3��Jͥ�n�wM�5qæ�6����U9���6�'��qO@%S�떱rx��G�@�8�9�Z����e�~���Q]�|r�<�f=ֱ��G���O;��,Q��r�b�nm!C��(裡�>�!qF��A��/b�)̾{@h�F@M2F�#� ����~�� �����^���t�	Ƞ���<�r	�S����A$R����G�q�̬/�u	��Y~�Np/;�ʼ�_{�G^N��� L/�,�me�H<��N��.��j���chy���"A����Y��+�&��7�T��F�����N��^8���Ʀ�x=w����P6�x �W�\᭎GYY����4��,��۞��PV�߻9^l�Ǳ� 8`��	���Vۚ�U�鷡o�E�m��'�3C\']&'��ׅЯ�]�%y��<^)m}�p�H���w�:��n��JҞ�=�	ƤM���n*ӿm.��VU�5�� �O{W�=\]�o$�y���䢆%T:L	.��D���ː�DĻ�&����>�;^�Q�Џ�n�O��!�0��Dm²a�#Z����I�=����A���hy�UoY�z\�i��j�����!w���]s�����b����k0��~r3s~`�G|.\̴Zh	%6B�x���{����rQAv��f&�b��d_��f��N!�Ka.*������YffH��U�+d�������Ռ{N��V��]'!������l&J}�+-T�*JJQ��+������yuų�L����E"3��@�Qv����'zE���؛@��c0P/�NN�Mz���i�KnI�rC^u���h�hc ɒ�d��h��ɝͮ�:�YQW�&�ߐ�郹���zz	�%�$�V���������D7(8���Œac���{�f�J=Ѓ!�$�m4n9���N����=�_�l}~z4R���� �u���諰�0�(�S2�5i��sa"w��*"%Fm/^?�0�7h�0�w��ν{�|�˼�Ӳ��p\آi�f`�=]�D}�j���_Ҫ\�ը7bG�w�C���#�\���	WD;��FZ�rBk~�n�����6B��m0�)�������E�e��Kw+�a|��:�& #mr�#����bׇs�OX�V��A�m^�ɶ*t�$P@E,E4�P�0BC�x6�9�����qfx8]YAHu~~�N�Y�EO�����ߌ'�!����943��T�ݐҩ�u{v�H�c�v=�j�;�k�b�/��=������'5�7��:I��H��H�O�(=ӻ�k���Ԫ��TCc�I����g��"�+)T�^��Z��I|ǒ��B�)�����}�;�QEr}u� ����lʾ�zn�;�x���� �cV���FW9o ��83���KYHY|�unnn\�%����2<�� �㭰�^?��Q1�(�)�;5�Ub���2���t��6���p�Nêj8{;��"��.j
���s�q��%p�=��((��Z�]jm A�}=y�0��zxO�Nw{7�����^������o*���sii)(Z�v{��5ۍ$����[ ��ʓ��;SJZ���8�����r�����xgp���p~��������*!�Z:�q/�Ԏ���|��=�d3�µs����M��u���qiX���f ,C�lK��[0�I�'���cw�nn~���H�ы�B���=�����?��H��6�4]+Ӌe	�M�I��8g���ˌ�<dq���H��W�v������} �KM:���<�s�]��edwt����G�x����@�A����%U���j�}U����F>�Lyij��/�ާ]����7��Gd�SrlG�Vy0���m'ά?��+ԍ�\�������7�6?���l���~z������Y�Ͼ���S-���r9y���!�Ո��տNMM���̠����1��P*3�C�7ZZ����x����UI�8+o���Q�IC��ҁ^�Gn���m��X��tm���u�eN�9���n��=/.��枯�i����o��D/T����MΞC�ZB�VkY��E���'a� 4q%�ȩ�.n�������q�O�E)��ڱ+ɡ�w��J�GO�ܫ�^��TΫ�ft�/����)���RC���Y�@
��o�VrC!&#�=U�@a���dz~�	�-��%��d�V��^.[ �G�A+Q޼�.{������т����͂Z>�iK�	�t"�7��y�X�w7��������OD}��ϣ��TI'�h����� DQYU5V�i\g�g��1�3SӔg��"1��XSK+������qٶWp7�1�>�cA	��љO06��������о
Xk�+w��:���`�~���Y-mᨕP���wV�n�Yd"�\?Lfp�D���Ѕ��0���ï�#/���E�Y�aŸ�v, �Fu���_�����.p���*V2��F�گ����P�uZakЦ0)�h����m�ބt�l,�UJK�����������.ӓ'b[թ�^Z뛋.?�+x+��$�n��	���#4f����C�3�(�@W�r��E���C!��Z�nnn���Y.;�tNvv?�U�З����9�O}Y�m[�C!�;�� !��s7�[HC�,�\4��>�o�/����L�
^���ߛB"������\�� ~#�l�7a�1�S�����E�!�|�[����t@z5���?H�U�j�K�OXT-�	ܹ{wy��k=;�	x�[0�yp��W��B���-��W�������?o�a1�����VB���|��@AK[��a���52M�&@}�LW�r�)vww?r�� %�wz����w\����
�ԇB�f�R#���1�+���$+��ח������ߋ^�P�Y�b�W��*}�ɴy�b���I��v P�ȯ��bjt�+�2*���%����
�"Ï1w�ClM�j�R�#gN	~N1��߿�Y�o�z�޼	�<|�AU�����,sN 8�.�S�C<z��}�� F��C����)�(��{�{�Wvl�ք���݀@l�60*�Hʤ����\TpW6 e��l=��^sQ�/iU�qi*ML����̷@98��(s����ؗ�q=�܄q�zQ�j�f#��(A�Ex3��x7T�>�ZZ2��T������S|�W
����B+�[�����[ ���C��3��ɜ�����, ��4pW �< ��>6��@e䍠�YX��H6v������_l�z�DS�=�C:X~1������;��؄e��RW+�\ɥ�i~�%�2�L������*�<�G�ڥ��{`Q �o^eк!|�uV�-�ϩ��c�����_��`{�g`�k0C�h ���:;:�e&=f ��݃�.�u���o?��o��Fﰳ0��$�Ke�wV������P� i��|��(����j�;::�X�=����!������v#���YB�U�y�< �h��r W|o���ASA��u��#n��9/#�:��-�u�� l�����p��[$�9�)ֺSQm���*hL���@�K�q_}�?�$�XX �F3��'Z�#ylS���͒�?���*/'�~0ձ���x]Ȳ<���������t�̭6�f^�(ˬ�U�.b�<̿��v��B�+[Q��qs�P��gh����U[ T���b��~���M����a��Zޡ�`�
q[I�T�u{�F��s�KHX�G�A?��Xl��8�H���@�@��l8e(���6p�	9=^$P��5�r,v��Z򯨚:e�k�[�;1��k��?D1�������EU9l����,%������m��=�vA��������������2+�Y��RRRX29�E������6�dA��Ϸ�]<��?��&z�[�p������	M�O�����y����	ޱ�'��4�mm}R�@Y�@O�h����`�d��S
8��6/6��8?���?+�K��������A<XZ���6�O�elIg'�>kyi(�М��,���s��g,�ڄ��يU�	��ZB��%o
1���.���)-"�$��E]�����	wj6ތ�=@(���nM�V쒮�:h[ټ�k���HyI���]��) n�eeeDtLL�@.��6�?"�;��+�;=t�����4�u;�P������{ǿ��M8e��id����}RzZ�8hpB�0*��f�N�����sK��xO����N@P`i-�nğ�۷�ʈ�0QL~~��[�T�@�EG;��X�^��OXJ{�hG��5�B���b�V.��-�B��3���\U������z'��Ѩ��WU�����	�'Sa��o�� ���c��v��T������F��۷o�ГZ�(�-n?v���7�,n����{;p�O���uo�mD�$ÿ�猧w!;~��`hH% <gZ+�e��߉>�:���^l�i�WUW���{\>'�����-@�Dฎh���Z𖖖�_���� �Co������C��x��9�����~v,����]Z0w��*��+�HG���t���HEmzA��!7�ђ�� R�gk
>��� �L]ѝ���ã�W�tc�D��<r���qE~��g�̬,)����N흺 ����!F�zO�[j)@�|Õ�o�{\8�|�/��:�}��/�A���)Z�����B�2i�Y�@��/�ݿ@�P��c��y|�;h[��FS]�,@�д�d`` ���m;v�Lpѻ+���Ddw��r������J�_<9�����RJE<���6�Ŭu��9gx�ā�_�7���8��i=:X4^���8ݭ:�N��>m���S�gŪj�X�S��\����o��'_߁w1)x���&x�O����]V]k9FBrS�揤T��}ӟEy���/�b��ZOe�RL��t�5I�:A�&���J�яc�l� �@I��!ݽ�,�{9�钤����m��\��\�U�];�?�����B�Z?�;�mԝo|���|����@�*߅_�,8�D�zu�2_�+f�x �B�+��8��ި%5О�1��D��m&_:;9���v��݊��v�����VZ���Ӄ[h��.���������wj�Ń��1Y�8/���#a&ae(r�t/I�5d0�N%�VX� ^�9o �1���-��K�b��S:��zݑ'�8���p�;��T�UqZ�+�J����e��a@��Q�M.�Xи��<�7	ԏ*Au3��q��sTqO� BT����7�����m��n�
X���d�Pk�I^|˨��IX��� N��2�z
�4=p_�O|I^����F���g��meX����O���|���%ѳ�^�'�a�X�˒0<�lh�G�U�������A�Bxq����wTQ��I����R������&Ea�Q`d
0-�� "|��s�Sp���}�g��U�
��� �蜯���ցѩ0����:�H�;�B#��`Č4'Wz����aA.3n�F |����ɟ��ў���ldH�O�7E�ΔŌ������'���3��&!�A7Nޅt���#�Go �G�v�<4*��|���������[�O}��ꩵݩ����%@a�o�?�Cv�*_b���ٛ9i[��+rQmgH��ZnR����z��v��^���������@��[p��2�&�{W�Bbp�ԣˁ;�lZ������e�d}����^Y8]_��OM��ֶ�mԏ�-����X
�@k���d�c�ù�A��&|��_$�����]<�c��_�K��eh�
����[9F�yh�vwd��Wy������Y�3A.��άVpG�9�C�n�����!y����3n��cTq1�-#j��@q�F(-��XM��'~s��=�\�Q�}<�~h���� �U�!�0��I�JJJ
�����<zI�y�m�gG���L��T�fiF(�{�@>�~�V�%K�����/�?ȱ�`�����}I��]����L�o�fz�&~q����������<5����>��C7�(�!c���O��Us��}lq#+n�����z�w��X\�=&N-��x�����!�����w�黄���N�����&�nz(x>�ؚ%����d?;*�P��,Y��(RҒ���3��5|��d`���v�y�f�P�/�z����� ��iΦ�1Ȁ>���@��c-�E[_�}o�����7���?��8?Z!��ne��P��b{t��=[�#N0����mЈ�<FC�s�!� �����x(D��~e�ڇ�i@˟-��BQ<���{]�Z��Z�tz��X��`�����5�N�!����k����l�PZ��#v�v�[U;ѕ�\to�TL����� |Ne5�L �-���Φ�|����G<���2x��͛��6��ʩLLLFv���� ���Q*��Q�ƍ�5�^���
J<�e]������Ɋη�`@o���$��;s�7V�#���fM��.*Վڎ��mP���K=Q�q1��c(���Ĕ�g��o����㟉�JK�����V�ldsiyPY���9�LSF�ao�qW�D��[0�5�����'�;m���N;�\�3����a
p|�ɝF��ƑN'���J�:O~��	�>���� �m�7�j;qn�6Kn�T��)x�Gzz�jځ�̘�����hPrN����>���>�|߀����y=��6�U��t=P��Z�L����  ���Ug�8�w��h�DF���P^Ss�/��ʸF�?��`oɗ��ŔC63��Hi� X\趻�]U5A\����#��� ����&+���p�EWw=zf� !��� �wzJqߝ�b��RK�x�s��$�=8���, |^G;����F7Kl"Y��p/���Â���؋��9��+����X"�7������p�4�T.&�����ֶs�n*b����q�Vm�S���J�1��@���W^�5�p?���1&:ڈt�7�5��wQ��Y�����|"ZNd� *5�Yg�^'�l@D�F��!����^^q�z�����>�Y|�_��
C�j=����c�V�����w+	7+�'��:���8F�%�z�a1���$�Y���zA�|M��t'�j�t��`7���O��U��`�	�տ-� z�-��22��Ad����ܦ�)/�[S'&4���5R��v�_V'~�����*����܀.t-LH�o3Q
ޓ૬�%"W`w��GS�d�]��ܴ���J���%�0u}�j�8B9��Lt9�|�g�&��k�;?^}1;�W�B�O�ȣ���U���{KB\�����ob|�k�9���><\��Fbc4�|���(�G���"�2<�==��<<Z�55g[���VR�.%�cc�Z[�����i���b,���1;�]�?L��y��[���S��UN�hz�S��.?�Ԭ������9@��`�xE�q���
ɖ6	��t���p^U�����N%:�R��[��?��p*�rigOT�-�?ɲ ~������Q�ѣ�-~�N��߿�v�q��E1�
-���c�A\��Υ�Oaa��?k�p��{r�
�

{���O4�����{�� ���d�k��*s�lb����g(����%�?��6�!��p�������h���DK�����W�m�Ը@�JFe��L��������yٛ�T��{���Gܛ�S�~��*)�BD�"�Hf%$SeΘ!�<;8��2e&dȘy*s�̳#�t̎�8�s������~����9�����׽�u�k�}��ڜ�3����%:�K�2W+2E��=绸��F}n!�u^��Ct�)��(>�4������j�;���\G����}Dv�P��������[���R�����b�c����fd�-'
�/�%����6����/��2ȇxJ�$%Ϝ�L�
z�����ɣ"��`hD:5��C�������f��K�X%�~��QO�1�Zg 
�]�줲j�H^(nHź�>���r�,r87�x�܈���� �@�����2S]ni&Ǝ�!=������͸r���w]a�Ū�1���*�ƽ�
�>ƚ�T��nZ�nv<������o�fs��bٝ��̻y���Ft��,P��Jo1�u���(-��e|�yz��F%�"���yޚٯ�yNɇB���DG:��V������R�4����-�4h�e�L���K���(����_|�;�tI������"���r�=�RK��+��r�j ��&�jo��<�^��BUK���p����K��h�w 5�[��/�jCCUv��jV��s�%t���`����.���+�tWTuM���)��3���/�r&_}R���Yf���13��|�`\��V�B㎫�>a���YA���q�*�|������dWwG�O�N�]	�CC�]�tt'	�pGv��#����N��Ʌ#�G�[ݳ�e|;��ޱ@�g2|���8�ꙧxk�"߈}�G+��H�u`z��u}�T��PƝv�f�s�CEPW
'�eU
�N�N���  �1����X45�>}AG=Ԥ�bh𡅈9��)ɸ��3�1/�s���J��>?��3��cY��n0
�|�Ӕ���AD
��.�p���i�"]ബ�(���ߌ*�5�n��K�m~,�`-H�:�索�";W�����H���M4�<�ۥ�5�p��h�z�[��la�qђ5�>�(�E>+**&)g��4_;Ln�<\e9" }�R'n�Ra�e'�ť-��b�8�p
�?�"�	�u��b�q��G����߼�}ℙ�BO�hf�L���-���De������^��{�����3q�ꎽ�t-tD>P��§��Q�K_���������<�t�%ߧ&8�D�=�2�Š�EO-NK�<槓)��SÑ7��I����ZZڍNN�+[<�����y�z�B��_y>9OGeiV��5Z�6��V�QO/?����\K�e!g��Z�?y�}1��{hҿEE�ZL���c�nAA赭�j...�����2T����e�F����"��a�6��c��T;G�|���ª<�8�co6�T���)^�:aI�5w�[@�g.~�I����jrC�1�>����c���vB�DP�2�D�s�>d.�#"��}���w����WcgȺ�����u�*�k�D\���Fr�ms���ؒk���,_#�!w�u]� J�do���ݹ�W'NA�g\c8��,'<�Xy���r �U�_�K	v��Q����9���\JNd%��sD����,`�����V�6cJ::�Ҝ��		O,ma���:�>���a�bq��`��c�?&���,�1�:������R�HJ��1jfT�.��
]W먳>�TT>yvut$@�z 8D�u6l��;�V鏟���_~���c���8��hD����D{< �?`���hj�H$�'��L'T�?���z����>I7SXo�x(^�X[��u�����\Ϻ�]�-�G�w�xG{��s<'����Ӥ9��E�[��F�b��-%Ŗ9��sҗ���"= L���r�w�-$���Q@r�h�BT]���>�-�iW�j�b���Ҋ�k{t2X����Pɚͯb��"��-.���������ǜ+����T����4���{��2RRp��S_����"�'����Cd%|��+^����~�:d��/�*���J�`��~����5{''3����$ʋ�HH�M<��CB[��,�2�зw���MV�Q��侶b������t��>�=9�!T��n ���yfP�S�_��h��/���{�R��J<(֦z~>� �|�~OM&x������}�셴oߞ�\��@YUg�Of�O�+*itp���]m��	J*r�+�,͜SN��ȫ������rM�[:V}N�)�F^�)��glxm ��#�~��\B/i����Ģ����H;iɐ��z?�*�+�29������B�?����6��/��v,YH]�&�[�V�h�rx�8�]L��m��q��%b�%���;�1��L�O���ğ���r�d���M=��FZ�)�d���O�<��Mo)b䉵�,��6�s8b(!�K2�r�3������x���lZff�{���A6��j�Ͽ�N6������7�þ��u������/իw��L���s��.��ȓ�i$u�:��D��x��+�� P��,+//���ց6��be�����r�r@=��Q���J�{[	a�M?E�P���N��*LO�b��o!2�-C$3�[���>Y��2���(.�m~E�0,�#�H5�ss��ʬH�S۾����7E%�y9z�U��wMw֦�O��}ԅ�����0e���J<
�~���f�ڙ/���^�=*�λ�=k�ͫ�f��O�협[�jB|����M�GѪ�,Mf�-��J$(w-�h,:�&^%.�	�jA4\Y��d��5�َ�������<�<R�n��r�@�9Ef
�m9t�)��"-U��xV�cץE�W$�>�O��$�Z���?��� T@
5_z���6MU�;��VVҺ�6���2�3Ivہ#&\��|	��I>�5QS`rQ�f���2ו������-�x���d�(�CC�S�١ۧ�8���	[�����/���~>A�]]Y�,j�]5��m����	�����ެ��/��m�?|E�^O����]a�g���Bq-�x�큗�
l�?9"'Xbb��b�����7�ʟ�*����RҼ�ZY݊�屬��㔝��5}��5M\SUAda´z�r��������1���J�������z�07S��Ǳ&�wC�Ԉ����� ���=��	xM����:.f�*+�����K�a�(HI��@;b�ި���Eq�w����2��b4z7�&��OJ�"`mx�hd�s�����ݜ`|s�\��& А���9�BM;�.�H����T
p��7����n"�F��<w��G�ڀ���q]��6'�9{6Kekc��ʷ��2�}���ss� �/�����eֶk�cgj��>w)�&#0��`:e@��/���r�m��B�2k>��T�焮7`�V7G��ͮx��MQ����`\|y�O�e��1̋�ƃ�k� �&�M�k�U�F�h�wL����R��M�����-��ALD�M�,� ��ّ������6v��f�UHl}�Ε	�������"��G�xVU�*נ1�H�^�R��J̜����6��U�q��"�|4�8����1��RT��OKc��x��Lyjr2���� p���,kP,%�b�m>��-*�3W*��L�Re/�%���s*�}��:|�~\���ܡ��5��Q�)pu���6P�d]% ��+*6�K�_q��L�ޏ5�{���R�䉿�OV��=�V]�a��Y��3u:z�_nj��G�x騫��A�'��-��3y�t�
��B����;þr���q����R���⭘���j���khg�Au����Igoob��[��18D��}�]<��;�j���d{�]��٘;G���K	LN��9��7@��A�_?������,�f���[�df�J����ػ���	O ���4�d�s�K�6�0�aK�^�(AW�v���LEOEd�l^T�ܣ���F����#[ϒ�]l~���p�;f��a+=�����_{7�Y�v*7��|�H���w*�J��	�t��AT���YV.в�_��������7���8�T:�<���MIOg�v�ޝ�<���dI�~B��"0ي��Zg����l�|�`��<���V�@�Mk���҄�o��ڥ��n(ڟf�opAN�vâ�Ѽ�N�O����ᗂc��؞]�s� b��U�^\����� 5��,��1%=��ɑ����gϞ��� �� )�癭������V@�&^���+*�__Ag�(�&�࠼N�\+���`pT�1����ģ9���/5�fWN@���HQ^>9�t�6�~��"���w�e3�E�{)U=IPcE�۠ڰ�����E�Dm��Ԍ�t�Ϝ��4~��^��l��o]V�d�99C��^D�@mK*G>&^^堠 �3]����z'��3s���Jzv5������>�sD�o�Ȕ�I�C�
JF�wu�S\�'CV�<+'>���|S`O�-�TDz_�ݤ��G�||I��c#��Y�IM(*X�/�"�گ���M��L�q*P5ۋ���
U��n�_T��Q���ls�������1�+�O�hRZ�EDFϔE���}K(��B&�8/z��}=����4 ��ѻ�s�K�r�xw�>k_�n���SK��j%����8* �Z�,Zi���O�=�+s�z�bd��]�bQ��"�Z�p��֖���)e����+;��K�*�/e�pi�/�bƼ��'���ʒV�I!��e�f:x�Ê�d���oqq�FREŞ0�����@P�g=��԰/A�L��wvg�rQe���J�����I�9"�:��$^'4��%��c�q%>XAnI��	BkԤ��8ӈ8{z�B�\H�{{��w6��,r������'���H�������W33��~�}y�v�1����8�M)Wl�Q��e���m���a���1w��,���ٹ��#�����v��=���u�(�_9vuz<�z��P*tt)�x����j�I����ɱJ7��v�4%{��i�N�QA�����:��
]g�߻�YF�����5�/����ЅǇ%��4�qi�E[DT7�C6��2ҹ�~���4f]Y�=m��A��|{��%�+�I	b�F/�����(��&��!5:n\H>FԻ�삋8)!��EO$����$�c�}�y��t�qz
E��7?��v���1�H�-�*����]�@"��^�;�'���������:9S�5���:|���7ei��׷>9v�0{���^6�rPN���`�&�]��[l�����ǻ�CRo�Z�	����Q��(}��Xt�:]J�z��mx:P����K���#{L��#����%�DEt������~M^�/�郢�&��8S��r�v��ߎ�&4#WMt$©�ut���\U����e:�46ӆmb5��X��]�Z����ʎ�&��I�GL��,�b��|Es3�c'��O���C�#2�GV�,�q�o��R��_��d6�W�F����s:�L�꾗F���)�X#
"�hÜb��F;E/���R|�3�_Eķ~�풠g��:�\�Y�璵F���Jx�"|�u�G�<K��1ǯ�U (�$�dfQ��"��^�^�ρn�mϮ��TŚ-����%�A�����w��E�n���:I�[BטYM�b�)O(��Tҥ�`��QỈ�KPh�	a����QP^��R��@E�f�Jy7���u�)n+`���Z���k&��_���lj��2�=s�f\�a�/GinS8�G㋀�V�.C##�I�i)nv
����I�'�q-t��׸{�ՓONX��	�+F͒�Y�Э$�򽒾|����~Ҥ�wƿ3��k�҄m@�]i������n}�R��
Ӭ�K��tQ�LVf�"�i��DN`s��:*
��bf�D`��x�W;�yM�z��O¡����r�}7sT�f��WR�`%ui"4�píL��l�7%|� �(+�� �&�|�>�fg�Q���*Ԏ~lV������	&	�Z�5WZ�S!���ǎ���+���&�e�P��U��w]�>��²0�J�j,Q8�/c=�P��1�5����5�����?�ϐ�'�@��.�EA#t�X�+����2}XXys���`q�}ZQA����_�4���=��~</��F�_Wb�J��x����Y���UA�)j\)p[��$49M�K��?nā�?�)l@Ke��(�rJ�@���	B���vT�1O�G��7��sK2��Lܶ��^�V�QgTTi�&I�,�m��o���,MҤ��t�;���?��,��?��U#(+J�8�;��۔�C=�{a�6�E,��:�B����.�!�*��X`������Cc1o��<]SK���X�r�=����@zQ�����u��[H��Q����r�����DW	���U���	�w�a��������̯�fT(:����e	_��y�x��7���)��t�{�&��X���_R�D��t�6`z>Q��NZ��QK�em�e����G�垟��;^p���F����n~�31m��()	%���?4�	}��M�����S���L²LPK���ZDc֪������EE�U#�ۛJ��`�)S�?��K}�X=�]�@�q���|���e��
�Cc�@�fXL1���gy��3MJO���^	���t6*K���Ʈ*i�	dy�bO�&X	1,�?���|?�_���zq{�bd5�͂�٩gV��/�b�|��qY�9�BS{bv:O����om
�<[`&-���\Gs�e/)>��4�0��!QJ>�PE�(�U2~�jë���T��;�aÇƷ�,�m�G�Ւ`������匃�d��z��ZyQ#w��c� e�,���8sn�X�7�j�����t���1�����wj�c9�����1`��铅?���E�xM�]F��:Q���=�� 0I^���$S�QI�S�uh�������hX���d@჎3_4۷p��zV���oqgst_����}N*zb&c��b�T��^�S��ue`>�p�!��`g�g���	�C�ׂ����y�~�R��vS]'��xLƣ��? �}�4�1Bu7�;=s1_���kT�jy�o\]�f���c�3�J�{�I����62��'h�+�		T}��?H�L?�\ژ��z�:V��c�SU�DJ���b���	�x�.�jf�!$E*�h]�jɖ��f�,z$\��;��R�O|N�y�(��N��J&��� ��Hc�U��!��{#K}���$���BQ�"}�	3��'|ˉ OZy?��&-q�-_��}�����
sG:�6���.08�� �8�����'�����_��\��L���d|��:����F�W@�>	}lKn�2�da/Z.�,x'���2�@��`���K�C&�=>������}�Q��Ϝ�c�e�+�$A6��z8�_H�kw�b�~�܊���9#��AG@�T�1��Ba��g��	�OQ+�P�h��L/!��%����:5�a[�{��aFB����!���3~�{� �E*��o����R�=�I����}R���������&�c2�KRլu�Z,Z��
�̑4��Q���&��w�w�	*����{74������/|����z�@�E�$�5c+�9��%�|�������΁ME�K�O�Uu�{;Eu���,���|�`k8��ٚ$Z"?!
����Ye�Z��i/�^��Mv��?�����E93���8���o�wA���S�*����I�4��vMԕ���F�r䳰����AX㝒�f��	Ep���4�5/��&�M��0+�=O��|3��}��ʻ>c������$fEI᳣(�S/�0�.���a�hw��Z|�\O��уԔ9��7���'ǀ?��|�7�?�}t�#4�ƈ��k</ �?�PR��Pe���Q���Oqߒ��Aݽ�����z��eLD͏Ͼ1ի�]k��Ի.���ɞ�Z�J��r�rW[���i�_˃�"pG���N/�O�J��?�7� �_G���;�T�+�X�(Ӯ�����Qr�E�ى���(��2����a��x��~9��6��f�2�	�᷏xzKA!�x���YիBy	�#����?��]��Ir>Cf�k������`�!�v���w;�.�7�V��a�g�W�=����f���]��80����+LS�Qqg��;����c���Ut)�B,qRY޵<Ӄ������z��*jOj�1�t�i��+� �ƌ�UbPG=4��T�H���-.t�"9y�j��i���T����oD���c#��(L�A����/�V�},+�ȼa��ʫ*V�ާzk}���;�;G��m�7P�~/~�i�˧(�Z��u�׾ާ�>w-�����#���.O�>X��JWm��^aPGP��\ ZTʲh���to�<p'?C�b�[2'��P��F�������S�8���u��^�r9.�1Z0���#2|b��۩�rY~z<J^j�_YTDz/V��}�u���?�B@�m�Us�&e4�:�-V�ǋ6j?;r���0]�1��N͊?7��Q��s�} K�����~-�_��1�(�mg���IVޝN���k�Y��#�j]���}T���GO$��n3���;1�us?��s'?�������Q���bO�[h�L$�������KУ�����}��аI=������hI�-�L��;$���H/䉣Aa!~��VG��L�7�{��?S6������ �sR]�����3���g�5��+�0�d�v�n�{R�Mju뚪�����	��]��
��-�H��i���&�u+D�u�[|�8��T/ݾ�rI�\=�!�,i�4�� g��������U*.d_ߵZ��L6�3�����O��N���<��D�h�k�W�;5D�d5�7L^�y�AA����=�C+�d�1#V�!�Yc�cb7����Ch��Uv�Y�?��V�'Be���#!ȥVᣅ+�y���+��#�d�VU\�nM{\\^�8V֟S%��h�=�Q42__j�����&��'֮��F�\v���c|\�b���N�Mp�s�J"M��jn�i�5�i�۵�oM�ۨ��$ljqs���?�O���5�np4��G+ׯ�9�\k��)P����݉_���~P��ű UAq��!�=��=
����Xogl9'=.t1(��S��K��Q�Uԃ89���X��R��m�%�^ǇF�Gڅ�7��B��`e��k�t�]��V�.S^T_flC��$�;Gu��|^�͖�Ot]��}[Z�	ټ������k6�w2�~{��ܝfb/�5�x��+�>���B��c��K՚]�6�(%�
��&���G�{
�m�Hx�����k UЪ��Ӄ�t�����6���(��߈����9�%����MSW���F���,Kok�D�a�ȁ(���8���"���ĿY����\I,Mf���0"���h���ٚmM�[~;�Ԃ��p�W���Y�����c�,y�5�3*7G�;4(�vהM�*;$����t���0��6:vR�����=�t¯
�$N�|~�=--�1>cغƄ���]ۧ���_��/:`�G����侧�H|�����A$&*B�+�}^�5��~�6���ZiѝO*+���m&��é5������I!q�'o1�)^S�BjK��.C*�{�0>�:����"�
.����G�|��� ;_�����V�
Z�x�q�66H��Nk�%9��wI�GS�]������R�mGq9���z�s*�mߨ��~{���9����R����Qe~L8�����K�ռ��T�F���n4d�2��=�L�����+[���F�;C�Ɠ5��h��<9��4�_�$��W���M���~:�U��h����ע#�5�W�%���YG��ZbEGc,��#�4�=R����|�� ��a��˭�Į�%N��H'.�T�RB����p�-�EI��+m��6-�_\���;gqU�r�H]������B�����8{ �`K1��1��rF�T��% ���+��Fd��Q�Ȳ��+8͖���2nIX�[���5P��68�8Gz#���S��YZ�C��-�����;�06�:D����/n\�����Ls9�!�h����"�vka���W%U�����n"�9�J�G�����RnN��W��u�zg
����@�����_��zX��8\�O�5�ً��F�5�#��v�0y``Y�4�|�N|ۓ+z��y��V��8���	~f�<��Q���vs�n�~V��i����
Y9������n9����H��߁�������K{���欈¿0���48N�{�`���5�����ZV���;����K�%�N�#���;-��Ñ�,���6+6<���*R(��I�\�+�ľcY� HX]hp2w���	�����4j���Hq�q�ZѦ�����d�����h�r��
�����_�\�F9Yo���-R ��C��6���fWL:���������0�%�Ytl��tK���G�⟡�r������@��[����/R^��ֹ� �J?���/)���2��Y/�*�Z3�'�� �b�6{m:+��n�VU���D2ʈS<�r|���S++ǩΐ3wS�����un+Ie���̯w!�|S��%Z�J���l���B�K�Q��su�8@��b,�)��^�f^! o}@��1�N\�I�-��o��T��]��=[9����"����l��3�XK��5'|)���������!��wPN��<&���?�]�-=D%]��P��4(K3wݝnZ-y%W����f�D��wk?���F.��K>{+��f>���?Y�t��]��w�=E!!L@#.�����k��M�<X�ĕR��F	�k�؋gi;/^b�l�4Y����W�<�fYk�e=�v�=y�f�`�R��S0��Z�g\��3�/s�#��?
�y�G<� �ʨ&��h�U������|M瑏��0o@��?X�s~'�7r�k��=����=(@���n�>=%�?�Wq����%
��E��+�N���r31� q%\l�@�d�,fr��&�$::�:[������Ī��8$~����m�}G�\(O������u�/�Q򂔬�j'�SUeZ)�oL��/���J1��n>`HYम~���=��g�U\�|�A�S�\�H�Lu=�*l��\�u;�
�+��*�)1����6η�)Ʌ�K�I)���r��Pݷ���n~�����g"�Q�Kt�d���\�Ԃ��F���a���5=��*��M%s/��9����'��Q5�*��Ψ�`�}>�j{.�{)�>�)����<�)-��;��	���I�FU�u�&&":�:V��H5�7g5���5��!�t��ֹW�)�pW&\%	���5U=y���v2Ee��JD ����SOy�V9�I�W�i 	�7��s�J>^�[ԑ��j��k5^6L!Ԩ���7�rE�`���=�t�!6�є����D���D��?�][Ҭ/]�`�i=�Q�ru�h�@���}��4P��D��S���W�[7R����X� EWY�G�`��yp�=-^�:j_�onF[�x7_  .��F��L�٦ƥ~��>��g�6T͇:������ez��t��vU��;��Y'��q�?dd����_U��'{$�������Җ�|G�"9����ʬ��S���I���(�OsY�k�z����rh�XP�z'}0ڝ����?J�U�[@ʬ����e'�ܵ�І��z����$P��nn�,��wN$q�xO&�\V5��E:R�l��	S�W>��M��s<0n*p�"!���4̹aR$��M.���f���j�x�NC�
<�;p������!��秪�$�nC�0tib���Bwo>��7�(�|K�J �U�{���HF�&j0l:�s�R�Ƣ�v-t���]���K����F���Βfz��w�U��E�Q�Q������Gyd�y�I̑4^�"%��%1�K��e靳��>��*A�#���/�[lY�C2>��o��54&�������Z'�𿚳++?��H����O�)N��O(	������俯B q���S��^�~�f6��p���V+�7o��}m�S��W�����{�,=9�[�t���?���^�{9f���t�(�3#<`-qyK]�
��&��!GCא���u�������r���Bccs�$L��¢��O�V�����C]o��	������u����%���n.5>�co僨�߫r�����	d�.�jjj�?��B��Sứ��|U䱱��ͬ��竸���W�KgMtg��`�n�`��%���rA�[�*QIK�����g��|i�uS
�'��M��������}c���s�kf�M�ݎ�zu��M����_	�u��ޒ�O���3�tۯG�Q�ҤYv_��7��h�uh`�����ɻ����Xy�G�߹J�$�t�QJ��WcY%�I�g��C�-oĸ\r��X-mw��,U�P�O�W�Z�۳!�06�{�	�<���t�^�Uka��B�e�������({~fNy���%�Q���L�|G4:X�̭�k��c���at���Er�X�QTQq�����V���>����&�� \$��.)�ŲPK_S%g��)�5<�I� ��@��]�UՊ���t��"�\.� }�y�~��%�:�fJ����k�w��Հ��^�	)�ݠ��
��N��.�L��yGM$�5?r�(&�~!99�}��)$� ��4&2��¿O��IE0ɸ�ẽ	Tl�����@
!n��;�
��ȷ�^v��|[��1�v��tV~`�Y-ˑE�u��+ $p��Mn����4������ѣ)۳R�� r��6��WLqt���Pk�?�k�\�����v!��@��ھ���{�E@��I���}	�,��ljɓP4�3�
|�{+?��1�FǠ�'�k��D�K�V+�����hK_�*�VW���۾%�>��X��l��lwc��1�bj}��:�V���P��ϻ��ߕS��5�*y�����U����3η�*�V��.��V�+χM��DVY�z0��±�t��h�Ū��������@�?�9pw�6;S��a�'��k�i욆>���J��G7��F�
����7t�D+���8����Q8v{-�:��;�ZM����1, t����["�9)�o0f�I�6��Z4{ԃ!������QաO��p�����+Y�qv��KY���O�� ��}5�.e���K��=R�S��)�x,���`��թ���w�1w|0�$���/�N#������S͞��K5.�шK�q��+�תˣ-�ntE�!���9���ى���֡��R��w-�C����5��8=V}�yx(�8�����i�!�=N�n)�y�?�oXt�Ym9������]���4ӯ`���ߪ�b��w�s*nY!d͏;��d����Y�\acg�BrY]��C��6e[zo��N�.��խ���[�џ 7�>{����f��Q������V,yCK�}!��ɐ�h��KM׹�ձ7dD K�/ܪ�[�7���$r�Lt��m��K��U��'}������H��Ը(n����A���,3+��U�G��[9��O�Ȧ�ˇ�ܘ�h\�át-,��"���5e�ЛFo
�n�ZG-eeeEY�^�GWl0�y+�O��З�ؠ?�l$8C.:G����§��99+�Lh� ��{��D~�e7*j�B!�b����>��.�%2���p�@�6~���z�2W� ��*�M�]X�]}0|��W~@�Od=���ʇK���翦���M���F죊�ׂJ�3��ǧ��w��A�w9{X[s�G�bp�\9��I��b��K����&�)w!s[�q��ջ�g����;������%o���W�`�FZ�#h X�Wۜ��XY��ˮڝ����Y5�3\}E�[{uJ#6?I�(�'�j���6{S:��|e8�0&�I{p�:���u�������� ������C`�4��Ϯ �����������ϗ���wl�[��&�*0-�D��'��<~�y��M`!�h��R���׳��w�-�L�]u�,�0�bt��t[��}����rh$�(JJJ~�6!�Hu�!���*���]���e9Gzz:j�9ǵ'c��c��e$�_/��?B�خ��h��O!�k��*�_��->�݉�X���ݛ�蠧a��s��`������T #��$�1Q���wJ�L��]��V�i���jױ�Kw�fш�a⡻��`�*p�_�yL1�{r�${�gbB�Z��ʗ��q�8��A$om;KO�iV�?\�`0�*��g��a{���Z>�U�ݩ��!�f���r�Ʀ�>�n�L��@yD�����ɵ%~#uK����3�q@4�� t��ޮ��6	{��z+�F��}��P9�H��N��E��/��>8���V�¯`@B�H+�$Ҭ7��׭�DDDz�4s��~e�J�UTUU�kח��.L����ː���:�?������! J���}6�6�Ч�}����d+ w��бm��12BO�j"d�hڇ=۫2��B�}����0�[VcP�CV�¤��u���r�ȱ8~�W���A�?~:��e�xLj�4�
]7�#�$l��:V����`�r���"0��X��V9�����L�� GVׅ�,_��&�k��P.(�jt/�n�&��'�c3�H�{�����6x#��r�1,�Q�ۓC4]�Q����S��@�Hڇ�����=�@A��e5�@z�$�m��*����k��V��n>Z�OKK�ɱ��f����ӱ3ϸ5l���g�:(@�������*LU�"��$���
B����*�owsm/�g%J�f�8�4$]�/R|�Ԁx~0�=p�$�i����kL!�&>a%�/B�[��pճA�����Ϊ�*$������LU7ʰ@���V�O�817��,^ n��!�R۩>�cc�n��̗��7��3��

��������d��w2�w�sr�]�Q ��|�;�&˛�}Uwu��g�0ǽ��IKM5
�������P�ݣ�5���0�Mf�/�,�T�����X�v5��Qt���!2"��q����(̊k�Q%�
��tS���S�l��6��EmѽʚR�Y�Ǻ����u �VX��*�:�Q���5� ��<�+�u<ؗ"�l>��,LZ���]�vs�H=�2����ǋ�r|B�{�Ъ�rꡟ&��zhU�Y�-�R[U3ڛ*�����{윒ZZ#j��&� ��CC[�I�"� ���p��dz���׭O��bf��F-1�w�D]bq��,�$5�Z
P{�y�>v��Y���-�ճ��&t�s^Խ �X����;&B�#�{�"~��M�
�ڀRw4��r��x�]��VŌp�/�s�K%'�ت��8S!�$4r͸"�Q�2�g&��Q���v�� ��qw0Ѵ���x�z�^������?#���ص�.c���l����+"	�s����L��{ҕ!����F��;,�nC)�Ɖ=?22r���������̥�˱����,��	�Z���Y�f�Iyf�I��Vi%j�.�U�(|
o��c;����(�bwڻ�5��Ow�ː�_�=�%7�v�.�0<�qͣ���B`d-J�B�i�n���>�g�x��5T��y*N/c��kF�XI*�Z�y�<GbM���Ę�0��O�>97�����C�&�m��=������l�.�8 ���X�>-�:���E?�����%+���Alv=Y��k0B��=��$]+�%HMY���ܻG)�	 }���*�añ�d��j��yYy��>{@����L2��4��ePg��x�@.�Ջ*���Nd��^�U��gs��ٛe�kܑ���'p�$1�Q��Pm2::�*	�4���q����\���� ZP�<��Р̏��⏊�������!��4,�c��|R��gr�vl_	��wg��U���(�f\�����bt�����^	N�|���H�*����_v^�&t��:������4�PpAw	$U���0{o��Y���/p~���H��L�I�v�؄���YC����O6�Hmnk[��X��*J�ޠA�q���w����>���g� 
p ����ʫ̭�	��&������7ՠ�'xb�+ў9ٌX�|��\tќv���g��Qߦ48�Q����Fh��w�����;�>������.R�	�x6�k⸶\��]F��W�5��&��t�r��xe��Ǫ64����;%�<�wN���+�����]���9:��\U<��� H*��E��5�-p�LJL���pv�I�к˩EӞ�n1�o����|Gb3���7�F�����t��������ݨ�Z7���vq���(�S5���֗c��K�pg!a������zʀ��-���t��/:��e���z2�/�T��0_�;�����h�4�n��F�#\��"�H���/O�$���ǽ|-�&�#d>����s��_���,���"��C�i:��[�/"��X[[�-��,���/K�7��VSgL�r8>8�\uNE[����9�[km&�~������x�Bk%3���m�Cz���{�_��y)(�:���Tn��N�e�z~EO�ֲ����w^0�����K-Q��X
m�?0t�A�ǂl�ׂ�+����1�I w��J0p_1--g�*��0煾���t���/a�c�!��A�PP~x-^畱�lNk��E����z��",���_�K�ʅz�+)��i�WlO�OQ90���p�e?Xx��X���S��-�-����#�-/�Rs�6���6:���V E�=&[Q���~'���+��\t�g�Ot���R��p�)�w8����ӧA��@���;pU�p^�5%N˭	�%���q\U�XJ8�+�]���(����0!$�yx��C���yW����a��;�A�I���A��6�T�V<�����o
�~l���-��b0��1�ښ������F�f�����%�0c���/�[G�lu_<�v=xz�~�Ťv��$��k���q2�*ЁR�TT��D���P�<���!(u]�ѫ]�z�{���ی!�Kb:�/&E4�}~�}�݄��&?:Qw�+;8�LYI鋃;�p�㡋��:yf�G���IdvA�q�w��u��u��N0�B:���*�������/�e'�@��<��K���mI���/%���oݽ�y��K+s��q�Y�c�Aax�^�Ͷ��1���at���t��3��̉ A1U� ��Y氰0-��x��t������)��s?�>�J��i��_���~�ڸ<�oaq�#8X��`��N����8��Y�!��
9s����TmGq�/W���.�Q�U��$)�N���l2��ܳ��թp�)������_a�� jخ�殹%5uԳ��	H��c�NW�9o,���|�*�TR\@$v�þU*�(Ɂ1]%6�e���݋�����:Jiii���p̂N�~ ?s�;j��^���K�i�-��o�
57��\<��)�%��.��_��*�=�<���� *�Ӯ�ҩ���W����]�Z�M��p;�v���7�8��,#]Q ��%���iX�^�^��V����>�?������/t����o�}"h����а8�DG��v愫�s�L��-2���b	���j�E���a��MQnK죧O��8��p�v�A}':����ލX^S�s}=˅�?�.;yϱ׫^hPG00^_J|H$}uE�Ag]�;sE jk�����e�x��P�qㆷ�W���ɩ��)�X��������L�I��?Ǝa�O=�SjN�[�|�>��(w�v�*�'���ů�_.�F�n{`�w �m���'@����Hx���ܟ��_6i�V�����!��0���P��8J����^B%��1$![�ݘ��}��*�(���Kֱ����b��X��}<_�������f�q=ι�u���u?�04,e�O$3e�H'���ԫ���m���ū���&j'���'�S�c�Ʀ?�+�b�x&�E~A�p"u/h�?G�? ��Fq�#��A�+C)z����s��o5)�����Ҥ&���?�����kbr�ί
[��r!^��i�J�Ud�}���1���M����]�
`�v�qu�J*Dd63�k8��?���� w
u�x���A�ʪ��R��$&|����/V�1p�u�L�	�o>\�o��|փ9DIvK��	����:����-�w?��iyT$:p��|UY�%��\�;���YP<#N�#֏:�X�M�xgM�x1�Q�E�G�e�6�i��ο�(΁����HBt�#�6U.��iR��ɱx;U�LKM
�Ҭױ�1m$�W8��X�ԓ�=����5��q��v6C��P�|���r���@>BP��VVv��w�	د���RW���:a1�`����s�%�eee�k��U%q��G�{g�-�bh:�L��U
�.��o�@�]���zZ*:@�dw�<�q<�wg��Zɞ��qI�������+��(�<���Uzl�as�T��� �1ۖ���s2�G������� ��eY}O�#���W�%�ŗ;t���O SZ��yy�$y�γS�+]"?��rI��8#�K�yjk �ښ�5k��߲��M�#��5�_�~j���n�x˼�=)�4���
0���j���z����#�W�~{�������N�Ǎ:_�
ުG�zz�|j�rFyHqc��/�QZ�Z_:g��8�4��a��r�I��=��!ʚ�ɳ���U��rr�V��K��Cp���j���?�ssv�z���6�ѽ^j�٪,-��U|� ���nk�0��dÛ��Z��tJ ��*�P��8�^�b�	א���"�w�h ����`&�TQ�	�/6�����i� �O��V;YBޥ�Q�D
2E�T�k�(Cq��6_�4��6�h�#P�����S�qN�$|	|TYq;���hz�����;���wK��t^ڕ�{��
<�%�H�,�Q�|e�7���ޕŝ*�+7���D�	�(tl�՗�������]�k�0�7h�\�ګ(�<�$Ek'�4͂eK�v���X���B'f޵�t���e��QJ���.0��^�$S�D�yW�O@�����43<��]��U�y|�	[�`�z�,3�	��ҍ����W�Yo��,��S�aQ�ߨ,nl�(7�1���D���0���p�n���
0��u�sO�n�l!���s�j��e�����lZ �������h�%���t� ������"L-�2��P�]�«�5�"�Q�� }��S�������[z~�C�|�ʔ8�Ay�o3k�/�y�#�o	�m��F�bEV���9!�
����D�Do�o����1��6a�k�O�&�{�j���q��j�~��^C����}�+���n�F���Jo��w�o}m��_h��-��LiE\0��8"%��y�ɢpRUY[�Jf�u@h	Z �iZ0ogT�k�5���X;f��	�� .��3$���k�nr���eA����]�{�f�s�c���R�7��'bD�x����C
��K[��!K,��7y�����R�'LT*Z�2�+�S��4��;gRJ�|jZKX�UQ�vC�7�}A��|#`^�O���F���� j��qa��;q)��Nq�傦F��#+�%�A#̖�3F��>�D�����l��a��+#s��mq	i7�x��>��>r0j��u�����͙��UZ�5'K���I>����j��m0e�������T�(n>�b����n�\�ͳ_�L�깐��*���@���L���KfLҲ�6rFN�R|��Ǐ��c~�X�����u��cS�n'kJ�i3J5}�9�t[�ruC���Ah�D,�������d�ac؟cqJnw+�9ڟ<�������`/
���3�U�${�&<�;����T�#9���䅙�qdh��;"�_�*L��.#����b(k�v7 ﺫ>��Wv�cmQ�/7��B�Bv�m��:�f���U[����>U��,AC�AG�g�%-�t�И�i)xZ"Z�oa���ԃ�Ps�,�`"�����Yc�l�hI�M=���0��)� ��3n�ѿ�l!ifP� �I�����|f������� ��-�i(h��Ìͯ��%�`�!4\[��'��6f"9TN�mP��X�t
�#�SS"��\wa; A
���qz�mlݞg(��DĞ�R�����3���ўb�,�V��6�:�{��6�Q��^���[ť�����!�7S5Oٿ�t�.66�?�N�X��wR� @ҡs>˨���n�
^�}���Mx���ՁF̀�w:��/,����k�kЮ�GJ�Q��<%�j�*<��F�⊶�@,;A�y����� nps� ��`�o�z�Npۙ��h��4�B���6�ZE�v^%�B�<���������zQ!�KP&X�~Ϭ_��
?�DFV�H =Ɏ	d�5�NGmx������ydz��������(��+U�`O����]�Z�*�����*�c���ZPg)��޺���{��%��V��K==9fw���V3�_��,--AGΤNL�"j��l �]cg���bC�҈�R�Z%!%�@��x+��s=�a]��� ��KC�ָ����@j*h���M���@�H�~ p�>�D&<�N�P��`�%G��V�n A>�hq�	���eqC0��e�GIz�Jy� \z�s ��LPc	9��9��6ut�$���Q*�e�!6�.�Z9�6]dt�]g��.y�( �_) �j��	���j4Q�n|Hh�kb�{�[i #ޙ�E�
�>��j<A���<�;�'SC$Ŝ+#���k�#�	���cuN���b)�,]4��R�_5�yt��#_�&�$Gg��J���������!��n+�L^��8۟�Ӿ��U=�(<��BX��Â�,G�h� ��+�P��.�8N%��cM{�|��/J�墮4�����4��6\�*3���/�`q�O +�	K`䋿и&��j�]҆!	�f�b�wݫ(yQ�9�H+{X1���)������Ax�ZN���RRR���w���(�MI\YS�|!�l!O���}Cj�/ �����Νϡ��'ԛ>F#�<dU��A��/�Y�#��T53̪�Z>]�Zʹ�\��[3Ӏ�V��5C[����Z��_��<��aj~�����'���4�]�B;���-��1�;h���+ s#0}q�h�θ[D&����]U%w�`�R�f��[�Z�y*Gн�xG<V6D��+��zcY�ed���g1�12 ��6�D�����R!�!pv\�z䚈���u^2��0:��4�|�+�������>#/�����;U{HWT�U��@��HH�:?)�)��{#��qg{���r��44>����	ʪ8���: kS�s(�{ƅ��Mv�y�ot�^A�a��kփv0,�t#I������2�����~�� �Q�|��@)��S�s�N�����@�8] C���]�ע	�.}Ȫu���ZI1!h�'�����ͥi$��YT�r)��� ��.�^3ؓ�Q���@|��S
���m-��\Ħ'z> b�q仦�"P �����Ll��qM�[:|��b~6��O㌍>�������"R<#&�B�=�T�f�!l�ԙ����1�\ps���|d�\]��L��B ���^e�|��m1�g�Z�3l"Qa�[XX�O�J��V
�τ� H��s��!9���u{�!ݤA�e�tl%d�^��	a8*ee�0��*U|�-���~��w%�G!��#ǃ��Y������ ��H�R0 �r����]C���lux���U�{}��	6����h����?#��Lq�d�@�܈�=�,{h'�y���t�u�s�9��
`,L�9�{y�X2>O5}��90�Z�.8.����[b�1��������>��k��z�iw66�6	ճz�~�02)�%p�z��]ͮ� ���`r*�_ki5��bdm�O����;���4�R�z uClW�̯@ns�rdG6�N�%x[ˢ7���5�Ri�5�.ѯ�y�E�H_Ej��;�wޟ�� s���,����j�@���.0rKC�G�^G�����q~@����1G��&'
��!�L��6��[���	�_�X������'r��I�I��wu�7K.�(����7�f쪩��;J���������9��Ug�����ӬgHGh�L_��W�=
"��!��+���`����\q���'k�� ��[�p/���9�kYL}�?�2�;T�y�`N��}j|tgVbs��x�3�0�3z!�����C?9�k%Q<��5[����5�b/2	���l��) 2��ƶ�='�ҳ��jզQ�����pN9���.�M����R0v`q���A�^Sj�_��b�: X�W�� u��Ac 1���v��h��d�Q�;���������-K�z���'n*c�U͟Vcȯ�埀�_���Muxc�e�t<����F$�q�n\�Kw������R��Y[�Y9((������x�����1;��6 9�v$H�� ��Зip�:��_�L�84����&��@����~�\H<���2q��I���&#?���؉��֍c��d-aC�}j�1�U6���b�gפ�`��W�ؼ"��V-�����U��e�|�a ����ֿ�{:�݉�Ѹ
��HAJ�ٙ�>�R����?T�Х�����&C@�4�w�o��k`�~���g��o`` ʱ�^��
�1E��m�M����<��茰5���*CGȤ�<��T+JM�	
ѐ�5���^Z���}���ҬA:�.����ؤ.�_o��8F����W�7A�F�}��?ʭ/3������9��Qy��p�B�۷o?T������̖�?ZB�F(���nV���<6��%1Fo����[��zf����Ż�|���c "(]1���Q"�q��%D�Rň:�lD�*}�-��e�Bv^ŃBi�0}{���t����B�6�e0J�9�y�o${��.xK+Z�tL�r�~*>�������<f�����5���PA�%�pƌ�6��2|�˩�f�c�**)-}�௦�`��8wnS�g���;Z�Y�a�d�+�Bw}�u^�1֖y,�����/M9�D��#K�����9( ��o��o��d����kg��`�@�9��¸�ƦY �p,���Be�'��	 �6,~u"4fS�ZM0�͡W@��D�"<?�4U�r@$9��:�6��P�q&X�Z{�bg�=b�t�<������LH�O��kT$�IM� �LS��k�T|M^x�'�����p���f��(5H� "%��+�_/E� �J/��F�n��� :?�]XQ������"�#�B�M5��8">Ȟ1
���>¹U����O�A@%d&��蹄�_��4`ۋ�`@�4Xo��a�YE�Kw���L�����(���)h��ٲ�R��][[�p�.��Q�
�_0rSo-#o��++p�����@�����Z!�Ǉ��~!�ƅ�x�	��~�AD  �:���9B�7�������r��%�8ޯ=f��XU�\+W~ �-�����@h��VG�S����+<N�u�����z�w`1�Ԙ�/$}x���ia^|4���zꓲ��r�ɒ��N�%�XM�bhs[�x�t�nq�}[/�%ϳ�J�� ��I��	L���vV2+���ܠ��?aܝ$-�Ǆؙ�6��/�Q2ҁ�c��O�Ϥ9��H:/��V�W�O\q���cf�7	�L��)Z��'ۣ�"k�uƽ{}j�ܡ���1eƺΏ�Pgj$)�q��x0e��Y��CE�Wz*b>R��+������qyƅ���ܒ�u�������ٚ$<��������x�̔ r#Y�R:�H�X�%��B��647�p_��_����	=� 8D�QUlXvD�M�g"�:�+M̊����͚ ���j�9x�D��W�/h~���ֻ�9�EU�"���v�Sk����J�>�Rr���U���%eۣ֩�����+�ĝ�|�
���N2���xG�k��� �J���ǣ!�Ѣ�bG��~~g�P3_�AG�y�؇$l�MCn�p~! HF ���&fRRR�.���J��U ��v��b8�j�a�#�|��L����QD��e&�ǂ����@FQ~�5`�L��"�?r��>a�q�� ��)��pDwK�t̮w+�'�Jf�L��ز��c �855����W��m�D�W�;��R�>��k���@T����6���A��j n��/��|.����-����ׁ��\ږ&�6��VD����l-�?H��{U�YIch8�D�J����`H4 �=�3/z7���A\ׇ��~��B@;���w�ݙ��Ț�d��2Lp�V��e��d����ip_�pI�kd$�U~�ڲ2 �Ux� �>��-LcP �= ߡ�Qz\YqAh~�/�Q��y,���p�eҨqibQB�����^�����v���3�6�{�d0���V��X���eѓ"r��1�er����^���+�G��rss�]����b�~ J�@�%��˗�ξ�L�����Rs:���Ho+��ܫ�� ���:񭺐T2چ_ҟ�^	T(�E�\��� cg��ܣ����BGO��O�Ƅ�j�m_�0t��HhOooإ�p��NO�O�F�-�s���gH��?��&��2��+�Kb�r]&��Xx�N�$�H�
�u|�_VW��T�ٮ�zIBxS���tõ���)�e�xQ���i��4x<v��a&�s�XArq�E��.��?�+X]�������^��p8��s�1�A�H�C���<J�#
n�C'2YM� �<�����C����\��I�̕��*�`Y��A�a�h��# ɼv�`*�:����zo�prZ���xڒ�S������5���YT<U��rƂuVv��.)ee��m�f8�`�u�煮�~�)II�{Y �O�k���L*�B7��{��쏯6��Q�U�_���h���� oKp8Xo���aa�b���;��	@��ڪ�� �۫���G�e �<2�گ��Ã<q�8 F�V�L�Bs���Xa�=$"{{� W��r&%��s�"�#P�q�Z���	���O*=�]�ཽ= ����<t�:`�ݵA�o�Z����WM,�'.����������O��ɾ�� �P���!u��Tൻ��e"���9�I{��E�*�')��y�M�/B��Kq���\,�_y#6�Z�� c�z@)԰Y,<Ȃ��~����(qWۭo3��V.c � HN�GǳY{����|p �)|z�"�{{䏹5�NA�Xb��.��	|������ED�����D��������U,�����I�[��!LS�E %4�y�{�d�5����A�~�3�Ɯ��%���<�~���|�S�^�sSD��mY>3�����s��?�T�C��x����4�%xIu����u�M�ˎ��M��tZ:�&�UU_��|ʄ�	��F���VI��$xW
1'<κ)|J�9O�Ç���/����`�7/��8��hvݯQ��U���Z��;tn!��-���6����ʜ)�e�֔���4�ɤ�@���٥�ƈ����GOp�{���s���i�"���Œ~<��T�M�K���QJl�te�u���Gnb(�<�ߝ�]ǟ�=n��A��4X_��p�C�E����
4����sU��;PMu�[������@�I�G�s�R��<�(������]�T��,�S�K��M��>�,1'//�l��Q���7���|:���}����,c����f��������=�\���f��~��T�� txi��D�0��+Ɵ��j�V\\�!Gْs�2�����K�ýsl�$K�b>���*-%�b����m����va��KQ��$P���m;	#>�'u[b>�l�A��`j�W���B �k:ҧہ���7�0+TK�{9�n��@��A�4���*�����w�T���y�ɴC�|�5�<O3�m�x��( n�B��'*)�_T����([�Y��NK$�d鼧䎞*U�|s$����SI�+t��C"��C�DJ������Y<�:O�6z3t{麇�͛p~c��������F�ա�����fB�9O�-h��!)��Z��X9�rG�zs6ǉ^��8����	�S[�>)��2�qGp*�o&��\	7�����n?I�8�3!�[)Xј�̴��3�-�����(��:�m�o�7y��kk��|�~�~;�+d\�%&fm�3�}�y:���z��I؜��=ٳ%bodR`]�q��3u Oa7����	|ܪx�=:�c6�[N�@h���Ն�^ �5���'�KD����)���v��ȵ��ӗ��!-l*;#�[U�3���`�"� �Y�)�ZVn��p��}u�3���qh"�z���z�D����ғ^/��٦A')Z�����`ٽ�֌�6�NX�h�m�x��vP�0����Mg
G4i	ߊ� �WN��֤:���8^YP���!�<�o���&���c�����;yl�+j�瞿�Ѹ8Iy	���v �OX�nܜi ��3KN�����<���R�fxG.�~�Hp�?�S?�T/�*�-)�5]p������u���X��9=����=z�f��N�=>捒�W.q����^�V�q>7E3�严[_����F�<���3w����f�&�#!\���&^�����8�s�r���[�'�6��(��ӕw������z��HR��#���̆�|QV������&�`+hH�Vo�����w�Q�@��\���a6ۀ��K79b��4S��x������ب�m:�Ҭt��|$y�u�'0F�D�)�5��$�	�묀�J��D�s��xC���\1zc��s�}v<Te��KvVA,�O
��/߻��+s�A��%����^�'��}˸�\{5�8��k`rܹd�ǽ*7��c�5���x�9�"Yn�����7�K������<ɻ=�< ����0��{� w�6g�[m�\�f��Z-e ��enx���qR<_zX P���q�{,�� ��	-80�F ��!2Ȭq=��w��~I��0�Q���8D�rt�j��%��鱱b��
zk�������8$3������V��?��3���J-�d�Y���������t�1�E]�R���(>G�*!sS��G�W�`�{I�s}cS���@�}���`f�I��_�-��P��*n���������k
ye�ծg_��T?�^b�ӌ�Ce�z�J(�i��V�>��a��	����h0�v�'ĠU\t&�*��i}qiZ���_E7�<LHd���n�b��z�Y[]�8�kⅎ\��c�,6���y6�v�1Z�9̇�F	̕�A�~�{Uє#�	����n�N���7�yW�c��3^�R/`�{1���A~Iuj�d-@�2�P�GR60_�'��!}� ���:"��(H�ߏk��H�L�G�������44f��7�Uj/Q�4����.�b��0�N/c��&Vr���(M����&׏A]IHm�C�	C�e��;bb���L)I�w��W��$�@�KʝׇIF���7��T���( �����v/��<�N���r�o/�\��,��b���hѢ�З,35��������Y{ �˹�����t�9w�j��_l~���P�]5R���	�-�*WT5��\�F򚐆�Nb�Tŗ���g���ܴbg�72u��a쮿��64L�ŭ���r^m���g <ݒ�h�'�x;;1Ţ�u��Ri#ێ�R3`�8�G�P�D�n5���K�Ldҽa��5_
^�$����S��T��������No>��R��,_�,�J��f\��pT��N%���U�U�'��wJE�K+H�I�����c dUw���@r�!�&��N�p��Sg�Eu|v� q��J���2�l����@�;����j�ۿ���á�ð^B��Ѽ�<���I�k�:T]��d^�����+M�pU��
�|�4�7~x��p4Vb�,u}<���q�0�����J\��GmG�}��� �ȯ�h���W�F*.�j��&j�HYuk)sn�� ��.<d�����:h)�1+O~z��zZ=����O���/ \�ٰ��8��p���LQ�5�*��$:�/��Tf����#r��Æ����qÆ���x�_�U��ЭѲ�!�����#�R=�C���o,]%�~�H�$epp0J�\�2�#�ϗo]��I}�茻6�K�4+/����r�cj˖��t��\�Z^��v�H�7��?��X�W2GV]���4�Ҫ~�U�2����-�����Ј������L�I���ބ�(Io������Q���v X��L<~�2�>O$y��U��;����n\��޻]>�����hIkS�;l+G�;G=N�@�����I�<n����H͒t��6�c�ylf��pr�A�җ�������`+q�/�ٶH�n��,���ĩR��xk�V�V���+!`����3��!Lm��'��'|�T�e�\-,������o�ߜ�G9��@C���aZ8-����H�OT<��ץ�)~-r%MO��;{/bO�[�8�i�=��Ro�zw�gJ�I�t�R����������m	��v^^G�F����l�n�7�PIܠz�&J�{��X�r��E��QH��: ��e�h��BjK�T+�*�m�����V���t�w�]��|�հ�a���͊.��l�⳽{��zθutt�wՃ�UX��WX��'u�����	P���i��M�N��J��Z?o����wÈIK�p��#F5��� _�ӛ`5>��v�������`�{���֑(lA��ױ�ʅ�~���%�"J�e}�bש��T���	����"�-<�dl��%�q55����-pn�8�^�o���,�^8�� 2�oދ���_+�Y.A��s�|ֆ2U:,v�G��m���ƍ���?�X��u\]�$�$����J]j�r��7���ɱ��e7���TC���ӎ����X�`s�R��ĿM�(�;���N��R��'�{QJ��Jj ���� �Tɓ��^>��Y�ޮ׆�u�N-�%"���ҩd�_�R<'�U�f� �_�X���&��;
3G�YC4���qII��n��u��ӱ-e�|�,;u,GW���( Ey����A&:�h������l.a�¹^�$���h�N��1�ӕ���{y���-�����7�^��/9��/��Gَ����P�xX�Ѹ��^��uъԄ�n�eॸ��}.^<�).Ԛ#�]i#q5�q4�4,���̠�	�~9~�sUQ�z�ᎄL��X&=~�ڑ���C?	)��[�~�o`��������[������ʅA�Z)��'���wq��\xW52wo�cܩOy��ؗ�����xVrF����&ڥ���V����urֿR��h�nDPV�ʅ<��V�v}g�h�v]�v�&�����n2�K%'��%��v*�fR�����k�>�D��n-�%�Om�N���;��ĜgE\<�����~��s�/]�}L4D��c{g�CzV���K��x֒���3���b��,�������$��7���q�wNO���,8�ѹ�%�m'/�i�ɇp�2
<tx����f�Z�t����>J>�aꊂ�hvV��߸�����6i�����L7ӎ5��_���b�l��.���4oy;�~MQ�_�N��uu�i�_�I
;z3����t�F�?�%zm(��K�IH�"O.:�9o�W&����Z��s��忬��KI��)b�!f䫹w�����cq���"\TN@c|��*��gݥ2Uf��L=S��+��_���	�Zm;}�����1�>N�nKT�`�w.g¸���I*��dϔ�	u{N�5�)�w^��
��$]ɼ�~��FШ��(�QӭA��9+�t��)�Wo*~�&)x��D�S���w�[1
��%gd�/�B;|ܽ�������Q!��ߑ1wK�lD�'O~�MO�[kiwɱ̛L���?�f?���e��Bycw��Q���X�4���Z/��6��K�����U�qQ_�;B�a��M�&�'C��֭D�;(�ðG��C!�-6b:o�f��R_�y�MT��.X�<������s*�@UW*��3��H_U��JT=���*nUW+���0�-u��r֞�r?���,oJ�+
��8���P�j<�8���w��ࠦ��ں���q�d'����g"�
�bL���:�_-ͨd�n�����"f�j����L?�z���/x��<��O񐚇!>�ә5ժ�L� �f�%cՌv{ۊъ��d"��h�B�d��.'=�*#���m��	$���j#ȟR۪>��Ш؝�-��I��um'��!��^�.�f���5��c���z@zY��M9Q�;�L�	���2���6���L�'���j^q���GW��$ӭ������7E��匐z���}�D<U�C���N�GVq��q�6n��Ǉ�����=�����{��6�Z�[����
���������}��'lw������a��~JW��3�w��q٫H3��ݡ�Ru����Uh���E{�V�[���V�><Ƥ�{\�4I[��B�38JG�w8�0���he��i�-��y��~���V����sU�׼f�Xz@�ͧCF���8�Z���D����و�
H(����{)%=��V��7e��0�ԏ�܊���.U|y�k_Pta�z<���Kz�,1�!�H��j�#�<�"˾�h �2��8z{vm�y��Rxl�vI���/��ijF�V�?�����yԐ�&������������	��"��Yŝߍn�����y��Z^��)�ܑV��V,�i]p��kk~����ϭך������Ą�̹=cd��l��uq�qJ�����Y��/貔�_,ؕ�	�uӊ�������4��;���KL��Gt���*y� v�?Ѓ�OW�k������l畒�V,�R�0��9�� .�}L��m��8����^��ب��N_b��+��>z���<�e�`AHf^�r�*S�����I.��f��i��@�96�>�~����W��U�����ԒQ�6��Pt�s�{4��i��/iy�C��!ym����D�絩2��'X_����EQ�Y	}�������	ܙ�NK�z����h�ׂ����I�MV=)�������=<���${��?׻Qk{��%��(�����w_�.��z��n��:R+�.Q4ܡ��#O%�U]�`���Bf==>�Ν�jfj��+^n���u���z����#�w�!�R}�Ȁ�94�L��������&7[�,:�I��s�w4����`%55�<)bZ��9�
jhh���ϢS���#��l�S��Uf��v?�Bb¸�v��S�/�
�R����-~�8�a�u^�s/�x�D季��
C����G�)[��$+��D"�t,6�c}I���c�2��}>>=SZ���6��9��v5o������J<��M�2.3���j���B�P� ��~eݕ A�vj$[�̕ڍ�u1�7�_S�������:�[�zw��9�]7y�{m�&%�_�Etr����Ƒo.V�hL��{��"y4�]��M3�bN�e���g���s#ͧ!�y)���D�����X�,F�%��'�Ž�&��`�@3��t=��Yߡ����l��+嚕Yw��M~��̘OD]�>�y���V�����p<`���f����R.��,�S�QK�����w*1���g~b�h��Ȩ~�����i�D�;r��r�~�M�m��ܩ����5�>̦��x5�->����z_�?��!��J��>','gV�c���(R�Z����׾Ԝ#�\H��]�=q\:��N�~ ��ݪ��U�x�H�f�߿���v���D��7�h���Уq���u�y9kY�+-s��!��Zt��]1P��L�D�(?as��Y�A�K�*�b�!-}x�[���үp���Ou��$a�e<&��K3
�qg���5��h" O��ΆR�9�gv'W�^����!]|��ލ��I;�Q�v4r��C�E�jLȩb}hY�v-t��5�F�_	��ߑ�3��[�f_G��{���
u��Rdil����G{Q���FbZil��q�R���a,O� �~<(�n��q=�6�Mp]x[8*�8� ΖX��41\{S�7~�N�ݳ�]��\
-� �+Ч37/�ewS)�V� &3q�m��df��_�I�Ɏ�;�d�v��B�7�"�䊙o��X�m�>=�?���aV�����4�j��[��0�Y4珛E���(8���w	P|[�=���w��D"����$�	J�槎����8�Y��j��gV��N�%;3���q����2YQ�nk���1]���XH*���͵z�.�q�S/��!���
��l��XNy��.� R�+V�+q�2s?��[qL�I]za����@�q�-�^_��12��.�D�E�FI��v����Z��42����P�������͎�Bŧ���I"͢��=�A����T��������~S����,5�2�w��oY�RU[l��cA�A�-� ޖ�C����pp���Ab�k���vv�毞��Єؿck��Nd�;�H|���#;�F�8О�EW<<��3���Њ�?�*6��O�so��tY�IM������X�TɰN�y�)��c��`. g���%t��AxPd��.�R
�g��(���܉�̦�҅7։��J���_���ԍ?k���܇�_���ߌ˝.�/�`��
�4�[�fKv!�*N�y4U_L���+�JY1<*�sO�%.��
s��k+��(�m����N"�V}� fI{�;�bG�c��lF���L�_��,���2��P)��DB�����24�e������	��pvY���,%W<i�����D������FI����;5�M�q>���'ڑ�k2Ŧrޔ3}(�w4C��@PL=�W���nw4�s4[������O'[*�oGz��ih� s��[�+-����#'3iפ�{�`��%2!\���ř�!���c��{0��)��q,�Eom��71��S��0��K\���ഒ��ߞƖ	�.פ�De�����^=�?E{�:�O�p�z�1�!]]ET6�_fz«G���Xab�J�͛W��SےI~$/�ܵ�ɐ�����^v㭿����eM�n3%���w7/,�oU�����j�f�͂�>���̅N���}·ⵢv�"|ӡE��k2&E�Ԯ,��>���O���3��b�ѧ�/�(_�8j�n��Y�� ݣxzs���Vm���L9�5*T�����<�a��x.ek���" ���A�n���hO<?�򼾻m9�;=ط��_�k���u�����5����z}pOb|����{�V���ʛS���Ӓ��Mz�xd��TCt�'�_�[�E.��l ���o�t]���Y�/��CG�1[��7�(�Q�~��z���yGb�6�e�p���&�8f(�ǹ_��}���uT{��V��VR��|)��Q+�~��c>��.��v�f����/ �k�^�l��	O~H���_͛�������i�`k�V+`�����Sr�#7n�ݚ�%RpM[�f�M��$Q��,�l�����7����se7[3Oca^�_~�O-�'��p���H$��ե��ݴ��젓<�	��B�u#_�
��"��g� ����^��>���:�� R2/�C��?��%�@��_��Mߧ��Q�H�<Y��*@����h=�-�6dh�}A� ��酭pH�u�t���2�lE�Dv�x~��|�}���W�>�䗫�i�N��͕(��� ��<rb����:��R��7��v/6�aG:VH¤!����o�8~omc�}��>B#ɣA�N�a��Mf
l:��g�����W�9"�(��}-��TP<�WY*K)ޅ���� �ݴ!��џޜ�t��ԝ��-��^���\H���{��4[Kp��*Fi�m&�=���ZW�b?S�be���pQ��O�z�kV�}Gڔ(�z�v�a?�&���$��œ�!&n��rJ����tڵ4~��jGܘ���Ǵr-W�?��#�gF���{C�����A=���EL�z����	"*�Xg�+V��3�!r�����E;��.�`���;
Ƌ�^�3j����l�\�`[W~���7 fz�2��
+gz�f��ϟU��`|c��#&*7�6�JZ#�b!����ޔ�A���Z)!g��3�2��L�Ft&$!�g=˫�VE;i���{D滸z̗H�O�=�)|����WB�R_��'1W�wB�ͅ8�.*]ћ�3����C@Zx�h���>�N�Ef�j��u�����������\�]�e���[O���\-��)��+�?���ߙ��,zW��B����aD)u�_�<-ӹlb��d������yׯ��n�
�8�x	�UXZ�o����?�A���5��Ko��Wf���ޢi��I�_����kZ�8�\_��ó���]�I�ׇ�������ۋS�{�1ЩA���bq�S�Yݺf����CB��A�����vF���=+��IJ� �q���c[�N�\�o'�o�JJ�v�j!?p���?ę�Ҳ��l�VgɃ&1�Z���ߑ�����4��9�Ĥc�H"�(�+��np˒o��|�"�D�`/����2ê.{B+��!�lJZL��������B�4�,Y�����ʫ�g�F��̠�8�#[f u�g{&�7���l�(�Ǣ;�f�)٬浺/� XF=oD�f�?��aW�H�t�g%�:�����,������k'튔3�w�� ǚ�D�`ƕ�X���S��_M`��,P�*�0���8W�[mjQ�4��\S��y� ������N��Sv���9�@&��,�"�ϰ����3b�����dV�J�Xut����A$��)vl|QNu({����~�*�t.v��v'eu�pKW��8�"��"ޣ��I!?�._�Y,I12�G6��;N��QFm�9^��]�e��wX�����{�P[�e�M�a��dřz��`٦+�0��.:��ݕj����X��;p��?�
e���g�K��ퟺ�!����&��f���N-19��U%E+���~gC��>��j�cO�fe�(/���q��ɓ�����$��H��X�+���`��� e���r[�an���<���k_�{�Q�s%P���k�,���W���az��Z�Hf�jYOz������~�/�=Z]�|Mܪ��'�(K�O*�(j;[n"�?��;�������R�UJ�ޣ(�&�.3Y�Ǧ��e�l�瑽�>�����}����}�����9�s���\����n$���� ����z'�����c3��	Xw:Y��Q��SvuU�t3�]�������7�i�/�5cY�tnnxg}9�`o��@����鐸���11�ܡ�gіW'�� (^4�}�c��}wAC}`ذF�Y}�����XN�H廭1��C/J��;�*϶s�i�^����F�d$��dqT��Yk�B�y��o XŌƕ:|�.�+`vN3�W��D���;3���qW���0���,�G8�:�o�,Vy���mL�OP<���_����_̓�!|3�^�~��N.� 5+��9-q���'�h�`�@�.�o.6f�{~��w�E��[����_|�6��';�M��!K�%5�3���W ���������d�P��<k��ځ|���hȅ&Sd�_�|V�i:���F�E�`㓫
�h@�9��g��hX�;���A�����	��/�������"7��蛪U�
R���6�ߟ�8]�v�{�ot��o"�e�g蹹�p;�
�u�<�x=�]�zHC����n�"��ɹ=Ʃ/V�X�so�b�޳W�>���t���g��8��!$���1��oMp����`�w0�.1�[p�E9��T�ǏK�x�k����4k�x�Ɇ������cO:�vs�T�t�D(�M��oJ#E���X���?��B~W�&���n�����|��orOkdj���?���W������H�$BP�jM�co�B<�)��P��P�#����sU�h�͜h�d��vt��k-�����Cp��0����}��е�q ���VN�)_�@����oN'
t[��C�uL}M�Ŀ�d���QI���n*�a}z-o���"f{�5 ����;;���*�7��?�
�I qM��������\ n5M3��e�'A��'����S��D�[𳹕�\�n�����
�y:�Kc�b�����r���������v�c����@|c�`lש��k����O�\W�|,)�၆-����ޢ����j����K�\�',��{��s�i<�3�O�|$�Ϫ�\�����σ��mP�0g�yl��=�������Pt�-�BWrgEU�5�xٻ"��Sᆕ.vV�TYc������1�/��w��mF����x���4��tY=����~�]��0V]�s�����q�'�����?�_�'R����	o�����������Su#������2���
/!@�,4>2�49�~g]���-+[���L����/^�m���񨀃+Awo邥aee���W�Zd�0Րt�� �"i�[�"K�<�:4S��E!��n\^����3�2A];��%�򕜻��d�� �߳��fJ�
�����X[�E6�n��&ٸh�֪E�d���F-�9U�-z_�\h�7"��F��h��8�eo�.!�A���w�A��������J���]�l�#�W#g���aѶ
��7��Ư�����ܮPB$�a�_�35=��$Cq{CA"fK���������L$��3��Lp妕@�-j�夥��x��[��N��>V�H�Ά�7�y����/��ly��tnmg>��/�`9]r:�/�4/�
+J����̤� G��I%J�U�E	q�Ә��)n���l�_� <泃�n/m F�C-7/�/��4b!B	T��y���um��Qk��B5�����K}O�;�q�2��xVV����nclѪa�WVx�Qs�e�u���ʓ,΋��|�_�-��&�4�C�|/5�t��E��p F��՚��q���i3e��qf���@�0*�5�]Z���p�eE����z&�Llrh��[�o�����)�UuN��Y�H�WP��՚�����k��U�ѐ������)o%+ӛ�������O������gmLM��#�Y};
�c�#��{N���<�jK�[�hZx ��q[`��­��:�#�]���!��¹)"q�v�M��~(�s�� %#�g��0B&��]m���ou�=a"^%�څ*;_���:w�,���Sވ�}�O<Á@�����|д�/���Aɜ֬la���C����V'�gb3�;B�@-�3�(D��զOX���鍯��d��i!M6�.����u�w��-`}�o�0%������(p���ԏp���zb�R�ȝ�Ԥ��M�������74�%� n	Tk�6��\�^M�����uޤ+�ZYXb	&3x��zE|��A�HB��H��F
{��f���z0Q��`��\�ұ�;��;Ʒ
����L�����CMq��ծ	6U�������0'de.�s0�����V|�u�	�8=��\nA��>?��S!j��{]Џ��i:LRO��dk��z|6�#�0eD�b%҃"��LX�	V������O�uZ�>v@�Pv-�Q���Ѵ�v�Z���K��{H��Dv��.m��ÆC��W(;�݅@x���սs����[&�JE���o��l�Y\d�mS�M��jP�Ðl���9�kg!7���}��u]las�D�АȻi�GP��Nq�=�uk�v�L*�ڏ�*ݚ���N�13�I�Z]�]��>+�f��~q���Oӥ`e���m!0d�bM���pw��ʜ����)[u�\��ʐ��`c���fM�m�G(m�rifm��m2��|6Nm�-\.��pYOpX�s��a��M��$��<w7�o`c�ށ�ZYһ燐���.��x=�5��#uM�
-.���!!��݊ A��r�1LAUQ_�G8�+T<ʷ��.������7�*��\*#I�
�����,MS"�	�jӲN8���w����%2U�oÁ`�x�66N�o B	U��T�D���&�Jr�ǒ�M�(�A�3��������y�O���XN��cᴑ��W�}��H��-`�E�mBW�ִGl�$\3�GŸ�ݱm���e|���ȁ��)����I�f;�!��Pq��8a���D� K��[�u����>.Hw�w�5R37�� Yh֟).��8[Zx;�I�F�/������=��t�j[�A�h����5T)F����� b�Vy��yB�:��H�^Y�����2泡Z�<������%]L���<9.�ݹ�c�o�=�����r�iA#�04s�g,?�Z?��7+y��7GB�]��/	��;��o�1�8���R����LYA�c� 9,Ldǌ��-�$�~(bux�_���J���o����+���w�c��+v*a�	�栔��0�i-�y:3_��}����e�����%�i�҅�-�CC�}�֦��.�}Dc��vpͼ�H�����uc�RD�����k���-2J�܃��y1#�D<�*�G#�i.JФ�1S�7k��e�ʮ�n��^L=�{1��lՄ2^��C�P�Y�2Όw�I4T��VuΏ��9�h�Xr�9?C2=������<�P~�rf�l�_YE�4���à�3�uWW����+�@ι⥒3m1��Hž��3�Ll�K�F{1f�M,"���� �%ov��IMNReg����ےAĆ�⚵��K�'K2�,7n>X��zYh��@v4�^0�Ð���?đ�o�Y[s�.�l�`6l54��n��ZǊ\%��t.���l�DHd=�Y4�	3'{:ۓb\�s�#�W�V$�i7�y�:z�4��_�Ѧ��H|7un�w�N��̡������B���)(ge�F�X�y���)]����O���#��iZ�D� '|�V��D��M!al�:�D�Ø�r�@>i�!�Kmmu7��E0��X�  �-K1rb����q�~��0����5��{�=�+�!��p$�e3/�|���~��NOlZN�#z��`�c��[_O�Y����2�L	���2�����۠���7tW9�7�'�x�w4a~��;E)��ވ����;?�T1�bO����dʓC��N�~Lم�3�__���Q�F-V�Ʌnr���'F�	�[H�DP����#ҧU�ޙ<v"c��o[��[�����˝�Ga����j�ǲU����y"�O��J�cdx�zb�Wܟ�"�m��bB��������+�Ϣ���;2�	��R�[v���yC��u����֬���x����,U~Y>U�0_s�8�i���gFk��]�ʘ����������T��\е��^`+�~��_��4��j��H,�E,olGk.��B�5���淃K,fF�k$���u�p�����*�5�-���r�Aw���d�J��D�7`�PM�l�!t��)G��
t}�U��"mGT�&Ʒ�� F����܀��BrrH=�]���d�5��k���>����چ\=#��aUC��S[o��j�\ S�-kWu�Eb�����,�G�)��_��}��q/�T�3�~C�⥎U|�ު�zDtzJp)���p]��?H�����J����Alc��}~/�cf��'�M�T�쟒����.''&j���QM_�����֘)&,iq�^ORe��
dM'�Tj�$Uџ��::CC����ŵ�Cg2�����΃����<y����fi�=�۾K��n�wz�?x��$w-u� Ջ��݁%c��u*�Z�ٝ!|�pO�²��l�ǔ�]O��f	��0�ש���Fk��=00�f�sg5��1?@D�,_k�T�Q�W��V��P�@���u�\��|L5w��u�C��0��[�����w���{O(1����!PB�⦋򉪖7<Y���9L*�6���̈́JVO�횛?.W�2Y�EAK���6O�g�O���H��a
s��0(������|����x��ך��"/E� �<���:D뇒T(j����ʚ�"K�z�1�r#{>)T�3�L,fd�n30ty'������g����2FV���ʵ3z�1>2��0LN���]͟c�T.I�l�	R�f�p���\_O�!���)�D,��BDg���O��(�h������K@V�+;/o���S�/5>����?�����Lc�Z~x^z�抰���=��Lc1���9?!�m��|�H#�-H3��{ç�@z����n��;���ʼ��e;C��c�*<�a��P����U���[���Έ����,N.�������lŗ ���DhY'��,KO��4c�ЈY@������2�bI�;�w�����6�i�W���_�E� �1����	'��kԉ������P'4$���`�}��o�h�a!��h�.v}�m�S����"�%to�Q{M�\���V��b�D�A�ϐ�393�*������Y��)�0�!��G��o/�t�ʤt��&���ުj\���5/�����˞,��1�<i�lY�y�bHQ�6޷�	,�=���Z�bk���'N���J7lۻ�q�4��өbVn�`�yT�4�&>Y��)�O����i���tǀ&�4>>VqflsB�p� �:���rޫ>d�1�ց��x7��"��'Y�~�c����x�JZa�IkL	1g�1���7��:1�gb�	�]x���v����e}XJ5z��-�
v����1�;BEE8��c���H�樦aV:K���^ZJ�n���]�Q4b���G�L�~$�6�$|���A5�ߘUj��ƹ~��-=����Je��c�|w	~����.�)�axW[
ղ/)& ã��=�C��Eoz�vJ��ó�U�5��W��~<SV+��PB#��34�dH��X\S�)����)���έ�oeC���ED��.e�.g�ʦ(ic��g�B��m�iwZZ'�py�*x�!Y���|}*>�i��7I�bgd��&��s���_��Ӳ�I���~�v�'���"�$�g�W�I{�曖w�О��e�,�.e��ӏ@��wj�/K��ʓF �"����<W��;@�qKp((�=�wf��% @��\zv��u&N��ְ�~B2�������ّ����*��ȕ�u����uw�]Q�=���P/�+�I��^�ѡ�'d<���/�/5�����|�u_�/������,�Nl�V�:�.�(W���dx95��x�|��z�Y�>��i8ҹ,�����m��g:��X�kU�}r��f�$dq�'�nQ0�zVN��> 5}}���6�r�R@{�O�wl`<���_v����=b�q�g lI��\C<�Aa�Y����6������d�/��eMKN�O˶�
7�Ȭ�۷�:���������W��VG�e�����HQ�@�UE��wiC��&�Jy��=��G􎑹MX^���"�ם���Ba̓�<�}���H��+0�3YOT~f��*na� �qy��Lo�k�M=�s�j
�]��n��B�E���z�b��9v�����u�.]#2����FA�3w��"���'����!Pon3ysP2�3ח^����6 288	��
�Z��`��Q�5��A���q���;�}�b؄w�٪Ŧٷ<A��4��kb�)7�<��L�2-���tabӻ�X��
�$�L�Y�/�����|Q{���wK�ʁٟ��Ypg�٪s˙{ƌ����F+��{�����P��Ż��f��֌&Y�xY�e�'Jk������m����(���f�k�@�E�"u�&t�z�����Z�|.����6}ʅi���� �?�д��++�"~!�\������Ж+"�n�\u���GP�����l�K��ޚ�yJL���m����8�pJ���Z/�hy�׶r�M�
��Z�
dсL��iBdn��?ɸY��g���-}�J�\�\�2]M�={���ܯ�	D�g�..��gK�q,T'^{�:dϒ2~�=5����~UV�a�K��i��)�2�[Y�X�ȁ=��oqfm³����j$0�j'�u����4�L��hsh�dȶ������ �����ۀ���|[ԷL��V��"b{�N��������4U���X����!C�Yn������'E������e��CDV�|Ȝ��pc&����O2�V��@ 7�Ĕ��]�S|,���ajT�?e�!A�"�9������Ja#�fd��F��}1ͼ"/�P4PZ�.B\2�*��D�F�N�j��h�����"/�?���+4Gd������
eQv�i��?_���M��@L�⒆�s����J́)�Ǹ�l%����f��Fi� �~4݀�[k]"8;=��_�<�C���䬨���E��Rt�XO�&��.�GF�Rb�]�u�,j�t��؇�|	EJ�Ki& H@y�ѧbJ���׭���Y�n�N�h���jݱ!���8��,Y�P�����-["n�iCp��Ш�%���R!������?v ��~nS��;.wNٿ�� �Hf �xR|TL�),l5���S#��RdsPWb����*}�%v�4�p�}ޥ2���p�c�f(ӆt5��kfg�vW3<l�1��-�a2�p ��,�J�V�ʤ���9<�|~�s����AW�蒼Y�ư&���a�;Xppz>�� �0I`\@wZ_ �}p�2�L}=��XQu�M� ��F�C��;���j9o>fR����B�ڤ��+�z�1��PT�@ �b�G��Nd}�<m�'>��e�����i��_�[,�0y	RJ�'ǽ=�yk�<��nQ�G$	�N���	e��%bw�*D�v�)lŴ���B��+��W�`�c+��4t_�X�ê0Y�e����z{��n�Tk��ؿu$��S�����g�m��>0�o"���޼�(��u�>�8�,bC��� TF��\ƪ��n�n�;,QZV�dM_0��ɨ�v�-a~n�zdZ�5����]߾5oګD��^3ۛ�'~r�������û��& �*(�4_@"������V�kb˕��颇{����{���cL`kf�<p8S����*]*��t;s~�е^1V��YOl��5��.�  ����^��3_:�Aq��|��.@��54@��鷔��V� h��~PG2D��պ{ss�߷|�}��A���̒�%�~5�2%��t���A��q�qЮIJ�0t�2`�@�-����j3�FO���o�g�T�s󠒞\B���Cz��sU���J�"e��,�ȢBQ�A�ۅg��� ��u�/��	a+mj0T4pp�_�*���~���-ԕ��E�'�	�c��������ީa�*)��n���`VJH6] aI�Yb��YY�V8�P�Z*�e>�ل����������z~3�N���>�e�;!�Ob&�;~ �Ľ�;��O:�z��La������Y���pє��+f�+Ë�@���)p�f�5?"
jᅲ��Jk�Y�� ��\I �g	��Ɍ�s;�fd�a�W�1A�4�`���
�A��yB�-)�G�i�x����k��� �,�D��7<��mo�Z���b� �膻�Zk"�1%&:a���*��4�_�)���i#��@-���7�:�[�8���:�פ�XVU��ws�=A�����載����Έ���}����,wZ�F�?��e3ռh�,}"Q�ElA�>`eē�K0b�k�2'�ʥc���(����#�c���k�*r1WR���2.ze��g�Ҵu����`��m��z�B�ܹ{��.}��~F���~5�~��\���5`�6q��0~��A�<)���wZG�b߅����}}c��Ŷ"�6*��L�P���i����`"�z�1���.8_v�+�:�:�Ѥd���/�g��l�3��j	Jؑ�o~�83f+���K�;�/:���p��"b��u���(���dT,��(o��y�Wq�����5<���xm��9��2[��x�����l=��;N�úӖ8�	>Y�}ZLx�H�t�=�Ά���F���]lP��j�bj��q齵��~���'�x:q���0+���L���������' z�	��^t������p�MO�2N֧�bg��cm��-���Y&���/��i�%�:X���&��YA�V��&���������*�j����in�~�J1ŋ��_������m��Z��'�,�� �lc�|���?���9�^8]�~{+���]���yNV�KhAGӣi��G������i���ƵUKӅ�G�<�����1�����y�&k6+��OVDٽG0�����{���⹨J�\'��5���Cb_�� ��ߊ�f35Q�d/��y#�s�in]�^i\�:=����Nq#�-�'�#�;��f�'���ԥö�U�w,�h�mw�c��GR��B.c�������K�ل��{a�����v�`&��)��cВ[���&��>�n˷�M>��v�E̳YW�m2��i�R�<w;�Vx�,�ϑ�	)_�g�Y;�[���Z�6H2H
�w@�p���Q__�MQ	^����d��B��c��<�;�{���}3�Im�Xt��g7g�}Ig��6�5k�]b�������u��=D�Zw7�W�����&%��j�	��"q%%����[dZv���.8}��k��Cg��\��G�2P�rI��d�������O��`�ϖbN�f���L����?�I�֓�^Z��jf��?:�9nk�.��Ln񴸡�`^��&�B��#^R��6wq�����9#��Ej�o%ߏ�&z�Јz����I+��{Gng���IaQT׽�fd���V~ie��h�kʓ�OW��dq���69�ݜ�m;#�U�2m��dj$��B�G(�_�H�J�|K݁,f�\����U\O�i��[cԮYE�!��
�l����B
c�xw>X��5������뾟XJ�TQ~G�Y����O���c`�1�a���Zb?�٩t�ٜ5�[��N�Y��F02=�6=+�"����FQJ�h��f8U;��9��V� �-�n��5�2����p=�À�Z����[�וL�Dʗ~e>�K���9i6��:ۉ�<ݰ��g�g�o���<�-��X&G�����<X��	҉*�?��L�	��yI�T�����_�@�4�]V�������i^�l�F��^�HH����6��/�l���c�H�xUА��=8��b�7�~$�MH. ����[���u��]��X��,yS��5��N���=y�-1H�5�2�4}g��E}6�jCep�OE�QVu���JH��4w�$�_9���4�k��D�iW.�5ѷ��7<���պ!����S.�N%���3����I雤�~����}���t��R�͌Ȋ�N1�O޳XN͡�9�	��'�)6S�����L��2�b/���PjxY�%c����>��V�]��+�`���T]=���?\�|�����|�<(_gQ8�cv���Xp'�J���v��<��͒k/Q�9�v���*��MH�q����L`���	$�Y�|�>�]3ܗ���;\��5z��@6��\,�JԴ�\���!��w?�XW> ��k��3-�yT�D>��8�-����~�(?צ�"+�©�L�>s']{a�Sqa5�ޗ!���z
�$i( ?�Q#��6�V8�Ў�/�S����&T@?���@��^w�kU�]�k�Ѳ2C�>�۳i�W7�8k��'�y�==jf��#����X'}8�7�l��R�f�i���1\�͖K�n��:}�Y3#� ����2�x~�-���-�1�O]�C��銽'�4)�@@�a��C�a�i/h�s�'C��v�7�F����u��GFBbeLq�8��Q�_Y����3M�r �欴`EM�Ar	s���MѷRIw|ӛ��	��jf�B�ɴ!� ��5���c����9 r5tɀn�)������17E�?��5��b�RS���Rf�YdfJq�<�q��_�J�?T~Օ�퐎�p�9�.dW	ǜ���e�^�EP>��i�nfS!|�´� ^��l��̄"s�
��m?�Ms�=�É��M38���|!�$�I@(�z�nJ'�1P�	Xv��z+-�T=/~�4�24ߏ�CV
� 6B���ϴ�%L�E��*a�6t���� k]�W��|$�^�q�$�v�Y�Hi3 �JGb�8�[���= �+{�.r{k]:5 �)9s���Ҿ�^�8Ĭ�R����]�		��)X0��\wX��P/�1=6�lz�Z�";�ϋ"�P��D쓼\�}�#B���T�OX�Ӥ�}�C"T! L�7�o�zM�U+���4�{�tO�w3�6��`<�ڰ�x�`c�{�m��ps�����r''���ݪ�+s�d�%d����L�&K7�8x#������nM�60d��cM(?x˸E��c��^���-x_�!��˝� ���i3�u2�Ht�L�oTtnX8��\Ƒɝ��Kg�������<���h�[o�ʊ{|� |�6&�"�����3��x34��Sw�M�x�3o�e����8]b��)���"���8��8���hKb>��:)0�H�#��x'MuuF��u�k�8<$+qu�
)6o�wZ�\s�Z���a$��n~"�i"�tI���O�XWj�?cY�M	qRLe�:`M�a����@�ʿL�M�e�a��IH��h�G��=(��.�,\��B4������)%�%Y�\�*�R�,0�K�@�៺�=�7ǐh������hs���ׅ�B�e���17m{�q�G��}c J��Yo�v蓳rY��1�����$�j)�}�H}�h#�.����83�^��jP�|��bf*�lFV�:oO���I�M����$!��l�0� ��<L�O�K�&�fu�l���s��l+�g�.��(��	g=�ɛ������g���ߚ�eKa�L��@�Z3��0NS/g� ow�p��Q@�U^���啈��Zd�u��g�y�*J�_�!����ާ $�q e�W��}q!�c1��������Hw��@F��ss�dy�>32}�`L��Z	p������� ̐���|�N����|�܋���HӰ���C��a~��cL��$�)�e�3����	�ה�;B������AS�7�
`ME�����D�aө�r[��k��s��벷���1��:#*\&�������@wg����{�A�lS ��n��mn��~U��`���k_���q�� R?��ږA��|���G���Jt]�"S���ґ�̋�H��J�:���׈���R_�]��KM���U���r���z�.�K����Q��I{�ʨ\#G~�3�{ɕ��I\�f�����"c%JℊRᇆt�_	u�]���tG��p�)�;���W�9T�]=b����>�܍�Zh�3��d��(��8��kÝK[�]aq�6�Cv;���S ���1�=�����Dp��VVX�%��A�й̹H����2�Z])�n=����դ����Y���� >�,�܊Z�.>�������D;����~s�h�%��̊<�kxb��4�9gU:���F����>���\V��t�B�e���Q���M��qj�o~6��	Ǯ�,o�!~&###�����4ɴ�*�� l����D�z �����x5��*��R��@f�I�~�Fl����W�`C2���q����5R���@�Ǫ�wC*�8 �MXrX�î�K?x�@|�U+��&�כ��Ŧ���Zݎ�i��`��j��ŉll��[izz��������H ���٤�FM���t�H��l�\�7--m�I{��nbWFp�Њ���gG�b�@ �k�" ���;����Ls΍�7(((���,�o�_ۡ&����������Ot֓��T�A i#�պn<��5P�2�C�%��Va�Z(�,����"}%���~UV
�wfՁ�i���|q�$�+|`n<��"�?�I{M��0Y�Ɋ�,�D�r��L����}���h�{�Vs˃	�[`;FR
�e�U��ݝ���ˡ��f1&$�(��/���(j��m��ȟ�������5q��i��,��"����+�iۡ/���+k%9���þ�u&s���2�`K���\Z�/Ǿts��GCi\w\)��|�Z�9�R�;�Q�Q�.�&ev��c�6n[��-���,�RaPEڢlSa��i�Y>`�'�piR��Ǿ�γ��w�t��=}���([$�X!sV�j3���Wg�$h��^;`�k7xn���x��vl·�Ǿ���0wY����Wf�r���`g�?�|�k	%%|�v?2�<1:
qe�0�C�BePP��
�����(~�Q��w�������
[���<���	_΋�{c7�}���T(�%�����ے�:�	�R��σ��$��ڢ�5 �W%�*�����-���m �V���y�U������0���� 2x��Ǭ�F,���oG�?���We�ls��ޙ�E�\�.K�u�*��YYY<B����`������<��b)������$O�zP��# rg>Q�B�d0���\����?��}���G�4�`C:��+ŧ��kBSX��ʈU��^�a6ik�?_��	�]�hb|��t؈��yF��������儂A�L����?����*!��|��R�x���/0��d���x��
���%}��9��y+1���g��y7�[�b{2��OE[�n �\Mtx�0�_zpwHQ��1bWr�hT���sg��W74�d�l��ru�ɳN�7N	P��h���N#E����&��'ǞE���^�������g�vh\����i|˖*���p���ӜR��]���� �|!�"o	e ����&73��k�`P�	_�)hin�K�n7�476�:&~\ߏ���p`�ad��պ���*��X��J�N�;����@ػ�,��r�6�� 6�\,��!g9��S�ee`�:�	��1���� |�K6��{�t�l�#�b�F���_$���~��E��J����dJO��IA6[���+72�'����v>>[ns���H}�;���|�Y��?3 �ѫDx\��ѲO�4I�#Vr��l:��Bf#ſ~��Z\\�d?n��۪P�ŏ�J&C�L�n"���'Z�A�'���@��ii��x��4�?P�T2����0�f���l�B���Jt�(*�a��/��q���k!���>#y:���� ��\{}|kyޏ��=H��8�⬵ ���\6:!xs'ҋ��K�2��h6w�}͋���:���6�UO�F�����!�2[S���QF<�u�=f����No��$%��E+ R���=�M�^��ր���.=����ҵ���]��sd�?~�cJNXr�p�pru��F��!: ��&���wV<����v'��Z����+-����_���X�$�9�k1l�r��ベ��]SU��s�R}r�
ZZ�K����O���^;ח������0=�ż��!�U	�xtR��{�vXW�^���� m�	g9��9|��ߧ�J�w@rv�Ͽ����L����O��Xb��G�_IIIڧЅ��'-J��V���10:J�ō�A�ӝ�j���ϳ�fhC���	;�� �wi�k`�
�0�l�.4���~)���P�[	�����d� �������a%��a�G���|6S5�����g�	�g	ȤϺO*� k"4g)?T	�)�?�t�qs����C���xR�1�M��R�L�~�spt�=��7�ivo�$3L�~U8Z��DV��D�tA����*T�OU� E�:"�#�|�N��o:��QΛC+r�rlo�?�]F��p2-{} ��/�xsM��	4{�F�3�t�}y�����&�>���=���H����-V�VC��T6��.#�gp��?�]�ܬ�p���
Ma7���a7���|���F(4+����Y:��u�]�f�[Lr|�9J�����vO7ӄK�{0�07~��	��:L[椇�H0������dG8���;�=N��	���4w�����nwV����o��ѫ�"�m�K�O���>/�qP���8����|��;�ԗ`2��&r"�δ���><�2>���;ߛ.7����2~�+"�w���*A�p��f�\�:��hf�<@n�P�>0�w
\�h�(�i�ԧ%d���7��U�u��Z�k�F���=����e��",�H?�Hȑ�9h��x�:o��eP�
�* �v��l�PB��rWf.Pii����ǳ��dWr���Z%��q��_}��c]G���is�S��l�0�(O�z�s+�0��P����!M���ASfb#����)n�=)T��s)$���g�Ko����PL}�]�B���6F�=uIs�]���#v����/-;�=e���@���ecOoV�*|cw�2O����M�i0\?�<~7����O�U��;�c0����d�+���p�}�łKJ��5�a)X����fh.]�tؓ\_�p @�y�"Fwog����>���O+T�^&�3���{S-�[���d���aޕ�k�;F��4"��cǽz!/����� ��E��yQqqI;�"����Fq�M�O�5�~e��sP��"<@}h�J
iGT���b2Ed�l%z�hcO>�YJi�-�`л7�a���:����6]	�� 7"�?�d���?BX����X|�\qQ�H�7���{�#�� ��?�_��NN����'B�^�K�V��d�� �Ч�#� Ml^��E�#��r��1�ϱ�̃D`��wv����5�2��r����[���[�ו'�m��~c��"뗞]ɯ���Mȳ��� ��s}���
aj�z|S��������ế���.��q��. �������Ldp���cGGǅ�r���5�g�l��Ύ@��c��>�b!YQ
z�'��79�@�{�0o�xw�I�z*����#iߛ�Y�ZZ�`� uw=@�xR;0��)%K{ܑ���>R�A�p�?*):�v�=���2����p=�'����׏;����������:���d׍
�OO������L�_���%��j�i�!�̜P��Dp'(�_��*j�t��Dc+���z���~�E_E��ֶ�`��
�~�Y�{�`���,G��I��ฏ_w6�`�ј�G�󢕘��=��Z����x<v�HV9�ؘE���;��bS�����t&F�#�c���~�`�g��agê�>+�(��Y1K�q-b����{���?%W�{�Q (aղ��
C��⏐�3b�`tp��� �]d���T/.����{�0r����5�c-�p$���U;X<�M�Z��;kj�ȴ��*��������/�q�
�OK�����&~F��[ru�w�����%.����x�ȆO��U�K���o�,XaD��v�}��<�geVΕl#N�p$H/V���c��޽;�#%'''lv P*�(��{�bܛa��G
`R��. V��;��+X9���K\1�g�����%Dv�p��2��^�����ZI�C՝��4�����<�(�@lˊ�=�첹U�����_��b�qK�������\������ʡ�/�Y �	���{�Gla��K�v�����]��q�����3�w���o|����A�A�y죏�ɦ�WC���6��e0��Ң�f���?O����J1�3���*c�fu����Fp"o>���"*�(pCs獾���ٸS-x9X%�Z���Cu��f�����\��W������+S��Z���AR,ޮ[��^���q�@Ri�*��1�Jh�;�̒�(_�i1��xNy�x�B�Bsʎ&�(ye�r�1�pq�x��"!>���%lؼt6yk�z3���/�~Am?Ȼ�ʱ�Y��qS��ībpa,��?R�f���n�ϟ&��z3%�{�hY��h�ɡ���@��"����v̓�Z_�����|&��uz�k���/���[�wz�Y�v��a��_�-�?\���
vh�e�2|�c��Gd�V 3/�T)��<L���g�8�<������,Z�Xs�ض(ɯ�~޴LAs��sa��nw�b.H����r<�t�8�ш˅���*���g��"m}`'�mԣ�7��sݩ��5ld�\��:q9) �~��w���oHb��&���4=�{��P��1G�V�C!b��U�������L��H2QB�E����WB���c.�_�����yd�Nc�$��u����W������|����������H?�RZ��n�Ö@��n������\�*;1��7���*�M��f�.��#7;Q:Q�����7��ʤW%x?�U�U�OQE���P�p�"r��}�\���d�9�J`n����2
�Y����R�#�����0δ�7��.Ǽ�K��$�2�F��]�Jj�vVz�sj3�7U���[ɒ�����o*���a8&��ә�B��r�P}CAh� xȃ������?Y~h��!s��^����훨�6�6�Ҷ��������1��\I��aP����SOU�Ƕ�jE���6�5���z@�GV��'�G���r��q/��;l�?�.�TZ� �h�Ko��.q���E��:[�Q�QPԖ 1t�S:uh:�Y��j%t���� ���E�h]6Z7_���4^<���4H�Bw''���Xd2����	��~�(!rO�32�,���'}K�$���z��nQD������������qˇҾ]��x�a����w+S�����߅Gmz��\�^z��þ�E���W0u����7L�Sb���#�ý20ެ�-t�}���#IBi�����$)�<���z�P� �kK�d@�j�H�&���f�x��h��	�@�uZ2�n�����]@[����1v xW�$�U��/��[��_6�	?�GS��?�-�o���	1�`�n:���>����J
!>h*~Y{X�n6��5t<?5����Ґ�9皢A�Yu��EVi�XX��ݚ�Zݴ�&���3�]�s����=i��a��~��%*IR2����������� [FZhز�c$�q������q%�t�y��uި~�����뾯���u��u��Fj¢d�yA�����������B�x���1���t��{�����ŝ�D����/�\����g�@@����M�m��r6q�%9�����N�!�{��dH�^.~n}��W˵]��9�Z^_�l���p'F�Ő֍^{����;��Ӕ�B��{�;s��,5Z�cި�Zma�[��͟�5y �3,��~M�z�Iػ�q�X�!fB�9;�_��c�Y��79�o �y����)x�a�U��Gj)oN���#����A}�CfO�kQAȋ˴���Old��"{��K��-�g~:~������C��?���L�n�Ǒ����H��8�/e{�kd��#�LX��V��BGPo�E�r���~�;�>+&�E�1<�wv��c���T���i@�~o�3v���vX��*1˫��ܞ����U����ugF� ��V���b�??CA��ܣ���ũ�,�o���H���-]��Е�MG�ޜ�������˥c���x{�=#_��W�~�F�`Q˯�������55zj��`��`-um	��ʟ�4�n��`ZJ%�Nz6f/���)&h�_�{{���&kmh��,ʳ�C��+�����-�'�#?��@��'�O,��Pv�\6#3Sa��k��5 �E(�=�ͤ了Da��`��`�����3��TuB�5��\�U�ۢ�Դ�4ҝ�<Om�qS�Ʋ^,�\�54cix��'7�@�-}�ۦI����F�?y���g�N())}�Ħ/cb�E������%B����4��՛����$m�V���_�
����&�9iO-��?�WĢ����D�(����9�RJIx� ��4�/�$�z�����L����9��K ֦ �G�,g���IY #����^�(�Wil"3Tsҍe��_ػ��J�S����ި��":��ѴUtv�˽�	�ݎ07�}Q*�v�{�g�6n6�|�j����3���[^s+ɯ��SvkJo�=�EFW��i���q�g�8|��=���`e,q�V�2�E{����$9+A%�p1�S~��cB#��0e���R���s����Z�E.�t���y��(!����e�v%y��T��<E�{�K��ؠ��+��q�:�tS���R'w���/���E�E��d>������x*^ұ���_�6���?s�G���j��C��6a�+c�vSa}�������S�g*+�Nu6����RsG�h�S�r
ø]��WF�f�t��$����@�7���P�m�=WL�{���<cؗ���t�N�L{���S6���}��܍��v�Q7��F	��ZG��9g��J�����E�|!#�k����U�$i��`
5��/1ۜ��W���V��*4�ŧ>�<�L�sa-�,͖T�*�� ӑ��/�N�����w:l��%����B:ؐ���^�^������9��a!�O�$w~N��K�qkڂ��w�J!n����K`έ��G��ح�{%g��½v7��~��('D��f�D�������~�=�gnԽ�*�L�i�k���~����3�|�@.�ѭ��SF���O����;�J������!�8�!����ȇ��E��n��w��ޚ%Vj.�FZ���m�H��x��An:1��lO����l�y�׷4�7c<A>ٴ�����Q�Nz����b�}�2Z����U���.�魊I�(8o�X��m��[<���W��\��ndq�(�)����6���#��S_?�2gg�D���L�ֵS-L�g�z	_`���]ߙ�謇�nC�ʡ28�v���
ʄ�|V6v�s |�������y��̄�~ϡ��
�����>�2�]1�q7��&Ħ���h�$��n-�0�8Ƿf}��X�2�����3LsY����\��`��i�P�+Xvg���A���e)E �Z��lI��T6��{�.ɼf�-���=p��/�%�
�E�S�{0��7�YK�~�/��LS����V77����%��}�`�$�p�o�5\4?$� !�����������P>�� 2���T����Ǉ��^�ū5��/�e������9~�忰��pvwYd<�����CK�8x<��&ɲ*�aT%`�.Ty1�V�ͱܧ�ͱ����*ؙ2��JbDV���B-|�zAK�tx�o�^xԌ�7�Q���/�F-���SY�5���ށ����	�mj'�ܐ��#����I�~�F��9q��:AfR��5�@�(&~���sϱ�\`�ѫ�x�Du���һ�M�7�^Jۭ�dy���MOpk�(t؛�R�1)���l��+C�zB~Y��X��5�?�Fk��k[N�wG������'�S���i��Hd{�Y�lo6�w9G���̋�kd4s��6��4��C���\�UM�O�� ��4���T�ٺ�)1�?Ջk6xid�ʪEw��%���G���Q��>�֪�4>P�f��T��.N(���]�n���L� �?�1���r��z�{s['�`�gꕡ�M&���4
�)C�#vW�=��N707z� N	Gy�\�gwH�<��,-hs���zfz��>Z�_���q��v��Ē�����bl����7
� ϧ�֔.�[q��Վ���фz���9�f|w�0h��y����v��C����;;;�3w6��99w)~�B����5���	crE���RD`I��Im�n7��P^q���w��wം,���)
�S�3V�ٟ��S=d���G���&�=x&�}��ٵ���1B�9�$o��jj�?'�{�$j�j����lm����!t�M�)~�ˑ�FF�f��x"�B�3y�ks�A���[&~��9����[%Y���d���Tn�F�|5�z��Ν�~�m��]�1#�UU��;s�%!2!���2ܞ���̾���"�2y02W�n��XA&S�f#m%aZG��.:��/��=�Յ722�Ē���5�n^�����]Yi����H�6�8�~�ŉ�
/S&�^�-q���3��@A�Gr�N�~|��?BΈL<�]=S�p$����c
!؀�ǗGH�7(	i��q4��Y~��D�sǛ�3����Q�	�#T-Y�'t����ݝ�\O�����;S"��!iQP�qR���x����9��H�}��e%�UpU���2�;Ro��E'�R\�w��\X��r�T������NII!N�1��Q�L!i������cT�7�\�>fĄ�}����3�����z$ �]X�k�dW.4�@�i��@e� ��s�q�|r�u����U.�w�[�t�@�Ϟ��8K9���BVg .(& ��|w�ĉKV��EX��DO�S��d��J�����ww/'ԯh��t�C1vt�H�??I]��r��y�G�&*��[���Рz��H���y��������@����	�kY$��k3��4+ �b<ՋT���@/�׬J��i1� �S��o��]�Thd�R+��[T�
��p&�EߎA�m�g��T����W�/�>�=|e�FS- 3�߇f���4����Wp��Ik�4��>L�ދmg�j�|��4��Uh�5���7P�H�$1�{{AFY������Fd��!��4B���G��x��rp�>��j��pc���p%f�d������~���/C��B[��s}}����:M������(����G.����Ղu�.�ne���W�w�5�S%~����3(:�`S��<��#w��ս�l	'_��y��'n�#���>����f���\����Pq]��nz���ӹ�ek�?;�7ԩ����y��7��޼ASQs�Ϟ'�A�$�O�S��ByXaa/���q!�*5�Й�����,��a�Y�E�D�xV�+���5ü�vR�	4��8{�@#�`���L6�\4�r�����N��fd�SO1co���
n-�icM[o��DûZl �(��dup�o�Ņ���N�.�p,�^��11‎��oMCV�����g��K\&/׸eʯ����c�7&(��������G0cJ�)L5���#|L}�a��Wts����u�F�u��3J��"��G|V�$��'��N����I}�V9��ں�LP͎�W�V���Sw�>���Z�N{<c���IG���Y�?S��3kO�����ϧ&�,,�F�6mt�
\��\虧�^J.Io�U7� ����Ӈ�Yc��p���j��թ��U1&��Y��	�Ǻ�k¼����Pn��6����q,N^�f���F4j�W����+Ob�;ͼۢL5��D�X�Z�o܏�cį�v6�Tg֪�$1>� ����]mm��&M�_�ް��t$�n����%%�Do1��^�9��U�qǍIJ3
�UH�T{�x+�`S��Y��sqT[E����7|�hulh�H6h���'��J�xV�V�����;�ɡGJH��N
�^�T4�G�Qd��W��g60�ljnnɶ�<xGq�����C��~�mN�y�W����v8 ��xS�
�oh������X�>�pǹ��L.W�ȹ��d:��5�0������wW[e��{���r9X������pU7����M��A$��"�`1���;srr��ӫo"�X���@^��N���[h"-����k�&H�o�b�uJ4>ϳnn���8�`|�apk��m����N�匯)/�+w��j����.rڹ�O���M=�v -���t�Q ���.זg��30Z���j�M���P�
G����ס!uv�<#��{�Ӊ�O�mx�;q�W;?���xe?���]١�1�zr_�b���ƅ%Dp'���������]�b�\���ܯǼ�M�*��W�fR��-��%���AK/�'Bf�0DS1��&�1�7���ԁn<�G#���V�)�`ة׽�& r�<Eў�S*�z��Ċ��B�|��W�
��z��7���2�XX��m�C,l���>�_�KM���Sc�B�>^.�M�e�?�Qw��[h=�_�	9����(P���(/*���O����Ү�K߾��o�sL<?8��=��d�e��q$�V!X��F��iD�9���G}��@{q`��WN�βM��<q����>�n�S�fCv1�����h-�E�Pق��6n9�r����L��I��ƕǷ�$�NSI��ic�o�^�I0���xo��A��E�����]�o%<c�̅G \*��Fܞ�<}�L��-"cfffʉ��m�x2]��o�S��4x��a��:�h9'�\>

�����t51d���[�3Ue}�)/�j�@\?���JeW�%�C�d�����u����Y䖲���w
�@�cnJ�{*#���kƆՔIخ1�[PE�S���n5��4�o�;���9nHZ�m'+�\�!�!U�KpdD�����;i�F�n��o�7y):����,,h���L�>=ɭ��V�<z��y��x��4np�w	j+u�ӥ��8�y�̩��#���]�<8�N��R�jk�]�I�չX"?��:o:�X@�P���A�Ny���>!����4K�'����,��R�ً��Y�N��}Z�4��M�h?�+�n�փ!�;�bd1�9Mہ��� -�

׾����V���#+ܗ���1J�tTV32�\�V})��X���KWWƴ�O׃!3�T}�L����a�E�_�"��m��6��7��\n�:
�ԩy/�Z�'���-��� ���`_�}]K1����>o;{��C'����RF�	���en�/Μ��s�;�z��g"�T_�B�(	��zD�͡���Ak+�`������
Ѿ>O��k��ȩO�a��\�1����A3��5�ߝa��j2�W��<xA�P9)za�	4��V�%�	t��t�[f--i��ik-F쟒(��9���[��:E�y��B�>����$�]��c��y]�9�	pؕG���1]���cj�-�zf¥��$���z�ɂ�I�� 3!k����h�~�|��1"��Ĳiق���G!��gfV���[p�$A=s��OfT�^AR	��/a�b4�8-�Y�թ�n�|Y��?��dk~���*q�\�T����f�5��l�
�\�4��0�J��Q�炯�Br���}3��>'E����A�(�7t�N�1g˾��y[^�F�&8-�>����s r�ivW>�y�guT��a�N�T�-J�Y?+w�S���< �=q��IO�����������jZ=��lfwyFΪ$o����a�n��م����\�l7&H?��s�e�W`�O�����������]>�R���g 	�����"�PӕR�3ŝ�k�I�GVT��x�%p��|f��j��X�����2��MUhJW���q{�9�:,v:K�ksC(�Ϲ
ۖL��ԩ�U�fƤ����6�kW�l�Ma�S̵y����/<|X���V���H���������0X֝�p�I�c#rk�a̛;8j���i2j��@ 
'�������V���hW���17���_���J����J5����������=EW��2_��M�*ͱz��.&���`L�~��E�y o�z�=��FJ,U����D�xͶ�]��pɌ���Y|�8�D�A���L	慯ֈ��&��t,�Y���8�>s���|^�w�Q�Z���)h�>$5� �&��|f(z�n�iz�(@��/���it�����tv���Y��t�[m�6Ѱ�#�_}2?%�a��i2nB��ABD>�h�x#�w��<�$�	��J��a�V���D��_%a���cQ����w�yLŊӲہ������S��R4�����=�Zo�U]<�`����a���فK�'���Ct+���B:����W��l;sAgqb�g��\���ջ�I��t��-q�ր#�srirT.,�hL���W��#�iL��ͥrv´�\�	\��ú���}H��Vo���u@����:1�%���l9�gD���YN�p��l��T��l]��ESk�j�N՟ ����7(�Jx?�Z.�q�dM��{�Bܢ���T	+)/���Ԕ���ui�D<N�D3�)��9;�?�8{�cR
؈.j��qU�$k�]Ⱥ�8*�t�0��p���l�0@r�R���0ӵK����Qn�[���'f�&��ɕ�O�]�ԣ��_�s J���"��lDk܅�2ӷ��OP�$��j�� R��}tѾ���[~���^�]��%�Q��|�*E&�u�L�r��� "p�261��.�'�z�c�v���L�r�zf^<poD���Pޞ���ǎ
FRV��s�p�'I�ps�����f�]����+z�ӹ{D������&�f�3�(`��k����.-��q�v�Q��n�2�;�~~���Z����M�w�K"=p^Z�W�~�I:�|�1�y�3��M�b<l3,�����oK/�� ����IK+w��H�%�������RK���+b��Q7��E<�yv����<��ڨ�/��-��ˏvl]7Ԯ�*� �IC��^���i���>n�ȋlG�-F��R.n��3��D
	��g
M�xQ7d�6�Q���Ʃ@2��4�64���W4��-2߰��Y��D\�@����3���ΌUY�]�!Ԫi-+�$~S��:���֩w?���r��o�}�0�L$�0��m��2'п����o/����q���N�S{�L�i��$��ߌ��QZƘ�/�^�nAB.x��ܨ���y�ĳe�S��&n����pgí���]z޹˙ܒ#����{�Ӂ��N$����"�!Wp'����+�����ÙJ�II����걕٘����{��m5�Y^S��
�~���u$��L�T�05?����
:me&�ڭ1 ��J��*�2Z��2�:A5�����d���t}M�F���U�-���zQ���8#LL;�����P����Ѫ�� B��%.�[�;�т՚���,�P�Qou�&�W�
,HV�z3-�m{�5 q�l����J�d��i�O�e�/+7m��GP�|:���G����to�i�YJA����7��>�1'������_�993� ��o�)4_���Əo��Q����98s��ݭ��e���k,��lB䛮\mu�&���F*S��O�F\���J9.p��a����G`���B��?#3��ԭ���6��Ni����3Id��X3������7ѭ�S=n��RU�}�;�y�OE:1�b���5q���a�r{�Y��D�<'����	ȶgR��[�o��KhvnU^2��v��/5~���;k_b���Y
TbiU7����()�h�o@&��o �L�ק��sXa8��ZV� ùb����g�jZ��dŽ���F�w[�.�
\�c�N��6�i.p���,�3�tx}*R@�������p�o5��sx�j���*�k�%�,���Gh�����-昑��Ƞ[M1�;x��A9�p3�����Wa���j���L?�o���B��Wg���ʅ�m�*ϡl����ˌ|�f,ϊ��� 4��v�h���'Tc?$�ޗ��#E}�r ��r�O�^9� �1<����YM��87d�_}"��Xu��X�͊섑���?z�)�C�g؏��gs�H��V0X1{)�盀W[���]��Y�����>���Q��@��~�O�tUw�w�ec���Q��m`:X߇� �� ��ΐ�}:��"V\�1���s>�0�T�菉��P~�(l�[�,��y'|�\��S1�{D��NYSFB��y��\��R��P�Rw�Lmv��ٛ{-{�dwl6�7԰R(5'*B�g�kҸ����\��IV��z����~������)y����O���ۨ������_I����a��~YT����!�p���ם��OO�>6��b=����\I�ҾbF 9�Z}�o0֏|��F�����#T��!\�׳�J}2�<pƗUзa�u��Eۃ�,X�]"��㌓��}��gau������A�X�c#]i�2܏d��W!���z��8�ۤ�fC���%/��gl�w�CS�-a�0���+.�8�u��+���|� �喘��fS��%K��[aǑ�Yț�JR_�c���PB��X'��5�m�s��*	�b@���Q�?u�}cn���t��?H�s��LT��nbSО���c���r��������*�{Bo5�/
���8=�7i5����i���!��a�,ḡ9������5rr�ǎ_=����0)d����NCUL�<�`��٪[N�⮶�#Y���'/+nC����� b�kr\pp�^��� v�g�g�執�'8�C�b*��٘�ڗ>��}'�&>�K
�E�S	R�MZ���_іhE�s�	���?�h|^�;.����X%BɉKs��wA7�[&�?��$���9Ch2���U� 8���Т�{/�~[��OS}�ȭ�=�wz���TÍ���v���ʼ2-��y�����2I�A������o�e?�lynܻ���m���E^��op�o�"Nb�o�s���&�Fa��D�w�v���苸�x�X2�bIb����֧>gf	Z�Wh��Ҷ���o�/�X
#,{�;�� P�"k��v�k��*�.�	*���V&����<*_�]4e�}���b�~;k"�f�I�A��;ݍu�%�ݴ�U%O����ռ�'d�M۫��^�v!MSn0�A_Xfc�M��_��<ae�3��V4t���{��2��eE�mwO���2����%AG����B�c�{6O��{sU^
��e�z�![�1��]g=:/0g_���u�q:$=\�ԙ��Z`/�޴��<��Vѵ?NI8u�)�G�}�e���>�ڠP�q|���ahp�<�!�5�v��y@a&��'�����֌��j��o0U����f�X��.<����r�yj>�tJ�o�T�F�J���.�_�m(�D�����0k]e�U��!�.N��z#���G�*Y��8�Ý��V{ ������SE����Ѣ{����Q�޼a�b<6�%N��:���ۙ���<+f��{��(��@�YP�*��������~���$)4���rȹ���H>w>�t1�C.�2���"�H�Z�� ��">A�kv�o��"�9��
<�;�sF8��v�Ikb��[g̩_SsA�ы,�dte��P�8bZ�٠��3۬S����#�����}�7����fWa�~���g�#�Ϧ�L0�ǯ���ժ���<k���r񮻰�S	��4�'_��]��W Lb!�n�|=���`3R�%����m��'�S�j��6=쉸�^ohv�[��yˈw��4�����3���ٱܟ��}:�!�3;��=;��H�_��k�b[���& \н��w^s�ks��T�}��ne����ρI5��1mʪOv�i`�p'h�
���0���;�e�l��*�CQi�/%�l`�ӇQ|�p��	���A�ʶ�٩��n>��/[���2��4�s�ن~�f��p��s-3��o�.GU?���_~3�x�)2T��+�/�F�	 �e����G�
�i�զd�EN����ѳ���F\ %���I1Ϲi�.:�}�4��j���ɇt�\�� �;&�ߛ�����b�;�H	�G��6������	�3��/S&��T�C����ryE��Y8Tq4I+�y5{і=�����qˍ�5P(8Y/j��*ݔ��]��y�|����R�N��x}�^�\�j���"�*��D���{x	�EM����x����ΈU��ܕo�-�N+����M�����+�1����P �:a���M���7�y_���h&b�jhTv����Q�Ş�)��4ރ�r�ُ��f�^��Z`�с�����[s/�z�,)'"=�A��o���F���#�x�cq�>��ם���j9�����
��U��#�R��tO�����)��^ש'd�ےW�e���i�V�j��  ���ȫ N�[��,Ugq�J��@����TY2�;6 ���U2�xpB�o��s��l��*����dTක��#����2�/�G�������v�8���6�ꇢM����
�ŧP�-�U�D�Q��,��#��A#ŗ�����
:�Ny�^�:����ӭ������%�5AoM��T�y]}��w�N}��3t�;j��2<�ȢF��M�4k,�����Fy?�"*�~�L!�=npk��P2�T�f3x�6^	��I�%�ⲭ+-���Պw?�7��<���Йߌf?��|�����o8��w�5Oȼ탸	�<!ϝe�ߡ*�NX `{à[�X1��H�)H��M�Se�Tt�#SH��9�5��d�G���A�ےޝf(��]�|F���M��{��}�~�N��F����lp��-���T�$��$x{{][%Q��d�e!U'>�%9G\6{���ڊT�� ������VUPt���	��p;��UB���s�.rZ��b�B�}+ݐ��X3�7d�g��9���l���@���8�v$%����I�)�E8e�ALt�hÔ>_ei�o�3�׫�R���!�AJ��cȆ/m�~���2���V���m��Q�ϚM�\�؊?���V)�4c"<b��Ϥ8��� �����!�T~H%e� 3�%b � |��.��uc7��U!CM7,?D&��O�� ���l�9`�=g(���f9�/d}�x�yh��-���GL�����RMӽ���W���O�ynF��ǝ�qi�
�{��y��V�/9ENn��>��t4P��b���9 ���ħS%�3����,����=N��k�*�}�@,5׭o��9��>|J����wAn/�Ҷu�_Z`+���{������wJ2���W:99a6h�n��jш#Rjў�K���y
��#I�ݮ�K����3�����؏�Jy��K)f��#N��m�| ���O��G-��׬�z� �	��8E�+�7͑���~�#.��鱉�#�eP?>rϳ���Xٿ�0Q������~򍀙��>**F���}2@.��G��������:;]�o�Ǟ`$;p'3p�0�!2���ƀ��S�V*�	�4���a�,c q
懳����緀*߃���/�$�!!����ipszꁾ�0��0��Ϲ8R� A�F!�Σg;?֖G��~���y�O��';1�[�0�Y�X�ݖ�fb��Ov����]=�1E�{���EEY�j�cD
��*R�=!<j���7 P4�A�>��*�b���;�W=-OG��U�]�d�y�ؒѐ�K�:�^�s��/����M�c��
�sؘ��ӴDT��r��D�㺧��0����Ŋ��Q���R��as|�1c�T��)���߂��WD���R���ՇF�ڑ]��9)&�G���g�=�ք����̩�pSN��� � ��HUT�Z }���� �a��W�#_(A�K��i�O�^�Λā��}��z�ϡd~�Ksݗ��]H-�-���ԣ�a���<�g*������<]�EɁks#��o!�U�����R���+ڞ0�չ�>[�+��O���gb���FT�)���959;�J����r��h��k����K?W��k��m�����Dk_"bfD,Y��N@E-�>j.��Q�����3�ɏ�	2�t���՚���!+!���+���] V�z���m��3b]��4ɍ �n2)� as�hƌ�f�?�O%��4?:Y���X�tW��F��h��%�Q8�h|]T�SY�i��F	�,���R�3��ڏ�JFJ�Sc�>��[|�g�vJ��\����u~�B��P)�y�%�WT�涚+�g�v���\�PU�������ǻ�h)~�k����A��d0~q���F��]�&7�`���y)�2���C\����?l��ʡ����JE����PC8���߆Km34tk�.Ѿ���B��E(R,N:W��ʈ_�fx_b�:���/Rw�
_�p#�6������r������rv2|lr��g ��w�oJ���ъ��Z�xH�.���8؋)���\�e�>U2b�cLJ�Ъ�z�F�V�9\_RѸ��U�-���@�H��[.9~�I��@�ލg�+(��f������!˻\q6s�����S�����ۇaHn�z�"e^�V4 �7�9#�Y%���cq4]e�K���7#!�9	��E���*�� �X*#�ٻ��<�K�<z����ș��5�;�Нu�Nv���	�W4o^�J��A�O�_f�}ks�v�G�+����
#Ŏ[�![�?�܄1ձ�ɦ���
�E'��u_G���P�[3QQ^�^�f��G��;��'�}f��X����(%V����1%ǟ�Fo)�鸌^6	�oA�X�g���I������N���C�x,���G�����c����G��=|��FȕZ�Q��=(�Į��#	8|E�t�W�t�Yƫ1�I�ږ"�kq�>�o�b41.)@1N���LM�rr�*�$�ƭ�������Jڎ~7��<�A�9��_	�N{ʑ#�;KQ� F�-�x��b����3�K�bvDe����/�����$��z�9�N�	�M�q@/��o$��
�Ο;r[S,��=�iS��|�/;P��t݈���}��!m䊮�����k��Ik����HcMP�f���-��M�7�L�W�Ƨ�����0r-4_#�)���8�4MX��~�]RR8�ݢ�>O0�h0��+�`UB
	�:��)ւ��1(�K�v4�GՆKsF6� Q��pȖ�w�Fh�P�Z�>�JRw�,Q�^�kQz�"lcҚ��s7�z3 ��憐yA�ڻ�V^��*��\��{�0'�N!���,�,�r���:B��H���&��q����'tW<`P'W���S�M�1��|�T���#jf�Q��{�T5x�7�����4�L���;��4JH�}BͯB@�A��mA()x!� ��B����OE�&�]x�]k�5_�׋���Ķ���T<�\��ȭJ��F��yqJ��wv�2t�o�����;��!E�������e|n��Us�����>Q��Kݣ�q�BX�����N;B�*&PO%�<����~�`g�Ｇ?��8�!c�> ��4ø&�)�ΞZpҼ2 }ȑ�����&.�[���3�D�'sv�x�%0�O0@ߙm��KܵTX'D�"W�k���$S���y��rZc�I������WɃ�]	uz��-3l��$��+
�F��-�2-�`p��yK�
���u�d̼�����PF\�o	�pj�t�	10�-����@�Pt����۬�	,yh�+��&�/gHg[A�>�7 ���c�XOZ�&wߏ��=��Uqk�Ï�����~}�gcc,.a�sL�m�����p��>v�����a 9<���ԋ��~�X�G�5Ov�Awޗ�g�N����]1;��HV!�E �K��ң�;D���
y{�*FA���ஂ�N_�U��~D��{�O�35�����dM��@i3�����h�������x�x@=��a^�Td��7���.Dď��ܒ����3[?T����Mڜ9Ts��:��	 �UOWi�x��
f�)�σVz�|RV{���6*�eAζ>pA_1��y��6�ʣ�A���Cg\n�:P��'ω�qzjC�(�O��O*��ah���I
�o��7*����Tk�>�x��2��7*E��� r'�v�К��ޣ�m�6�_>�}t_�On��w�=3[H?K.����
�Vn�ݲi`Wj�2x�A{UH���������x��%z�S�ŋ�\\B������`\7�	#'�<������IqW�W��.�1>��A_E��� �0�� b�M�M�R��4rN�g�)�p���ɢ�I<Q]��õ�L�J��Ez=������dlҰ';F�Yr�kj.)�6��V֓��"���O�o��7������{9�PE�����h����͠F�d+��Ĵ���OQ�ӽ{���`q���?M0"+Aީ��)�~i���G�C��P�M:fO��țz�D�G����@�R��`�A�Q#��q�����v6:�4T�Fs��{�6��sO�1)����
�`>	�%�A�����5My��E˅�Ŗ�ị~O�R-�����[�Q��ď�z{��7��CK <��5Ѩvɣ{��c�����,gU�6�B8���5�R�UN>��|~H�n�ܹ	��|�Y���{���ɯ>�j�RvWM"@2�+#[�^ _��;����"����c下}�C�������8m�c��:|n"�\���T@g���&�Yn�{��dTJܸn)�'�� ��^T���\$�����������&�SS�"���w_ge^�o�J���|��ى�D��g�T�\���R*o�
��>=q_g�c�ǆ�߱;�rW�	�L��ݸ[u͵�����	A����u�]黌/%�+�T4��\�g�<0��Ȩp���b�I��R�3eߍ��l-Q�[���|e+����X�
얇��fSĭK�<-�!Y����$���{x�]��!����T!�GwB'E��㹐�����=�Π��v�D�Z٠��>���,�
�Ôw��e!�R�Ğ�ݩ+l3��q�Eo�Q�8��t�Y�/��K�`Vq&�~Ա*�v��ƕ����M^q��4���pXմJQJ��E�;`�ŝ�Q����U}v�KJ,�mZZ���$݇v7��CS�� ��!|���f�����7[��R�_�2�Óٙ;[p+a�ރg)*��6��>kl�Ãs�;+�Fs&��gw��Y�kEÜ�W:�ko�ި���VQ0~���������G}�I⮈e�,��5)Vf!�!���ج,xo����HE>E؟.�KV��4��$�<Z����Pt���~G�_�f��HQ'�\��F��[�4>x|r�m�yY��h�K�iбS�9�4@����J�qt��s�[����*�/As/ _������q[CReK���W�AY�n�t��Q��Z?�k���+���LO�r����;m��y�ͮ�Fp���ĝ��G	N>�8H���� �A(T~-D���6��9^��0����&Ɀz��,�V�y�EhRᱠN	�l�?�1�
�$��ϝ��WD5�X��t�������b�	'>wRu�����*ϳ��s�s5��b�3��6�+���Ż�����f�G�	�܆��mo�DL�ef�%���V�g\T�S��`�r]Q��v�z�|��p|E�3~�Z�?>.�c�|�}���P;xƊ��4���u��J�ܸx-ޗoܝ�%#��%�6�h���_:�,�,+뎐������DOͤJ<<<��+�bAۏ��e���+�����jy!��\5���yZn��㴲S�{89��Ep%U�b �~��ɑ��!��w[�/���"P��2<��!h�5��	�����]+=�����ӷJ֌S�w7�= M�zO��Q���6�]~�\l�(�ؿF�3Q�5�7��"��Y̷9� ��O����%�[O�y|�)*)aF`�%�"��].��~��d)״ӈ����Onp��ð�o 7%K{�����?a���U
�8[�~��^z/��V���t�J��3;�z�5�b��8�¼<�LOi6z�7څU�V-��x8�SB�͙k���IY��r�(ix�������)PC�5�s�(ϲM�S%]���p`�fH��-C�+�\�N��/�M'����{��dC�Isy)��h�9���m���q�������_�w��g-lw���ٙ,��T9�57I�n>٩TKQ1�Gt�*ߙ(�HMM���4^�0�A���1����Y�%%��r���ce�y�A��ka�H�]��s�
�ۆzƔ�®�\3��H���G����K�2����d��q�k(*R���Tl��,@Gl���fV6��B����w�?��X�]��6�}�C�vW�����e₮R��ki���
��V�!|]Ӆ\�����\�MT!�6Dn]��������q�)))%�Z?�$�P�։n[-ϙ$�ظ������"%&���oLadd$Y�)R���O��oo��}}} ����&�ڈ6<c�?����C�rN�������o��QƖ��4�L��J���ar�GK�ꆊ��X6�H��7�|��^DG�+s�q������a栎��4�7�25��RR�gSݚi���`�FF�__�8}�6.���7_�K��NNg�W���Q�_MX�?��<����Q�DE�BBʞB��;!{�쌭"E��k�/c�cW$���m���������޿�������{��<ι�ܫ�R���D*���qS�%��P�����Y\\��vDSO��q�[?۬=��B�Yכ&��9L�1N����V��?�ݢ�Dt��Z�K�A<u���5j��]��+*.g���>|8�eT7nͺZ|:Ed��1���#�Z ���m�"��7I��cL�{��)�g��� Ĭ��*��I���|�a*�9\fC�$�[fϭ��L����w>ƨ��KH������B���pw������
;����_���-.�*u����Z��FYC��G��ny����i�4�������_!<f�[�t�wߚS�PI@�]1��V�E���}�]PnR �����z��W��ƞ�gѩ�1���~(����d��S��^�	,7��Rr�l6�� ��5_�`�j�ŧ]n�wˋ��P�j&�+��賈���RS��xn��4�长V�������4����c�;V����+�<`��{�
��e�Ӓ����^�+El2�U�����7�XW�9P��?zC�S���~����7����8
�%� �/�.ë�BO�����+��,'O�a1:*l�8~Y��{�zŁ��o����ΏEr��$�z��0ع�K����A������qp�0R���ȴ�:^��b�D�'�g�\�>Ө+�������5��`���U-���;Fi
��hA��*+�ty׳�#��n�S��Jq�]�_1��zh�
�9�������k�5ڏ����E���>k_B�e3�Fv��Qt���غ�$��떤�ڔX�Y}9�"e'�l�H�>�C�i�:�ܝ�:D⿃�H�ԍ��Y����Ik����n�QZ�P�q���.��'�G��)5ɗc��jSz������mU�DZ�@�.Uə;��S/�ƍV������*.�
1bT�����4#�M�%��)�����ȝ���sVõ���Kr�ӐmK�	���!����P���>��X�������	�1I����%�I��ť��*{��k߈��L*�Ĕ�y�������=
wG�R�-mkf�w�]K�4[�Cd�4-1l�V���*B���I���Y�{�u���;y)�h�t�Aii�����@�4h����kR,i�ֱ�},#�4��P*��#�9a�"v�����4����>c����@,��"mt�^.D���9��)�Yz9�=�@�3ߗ�X���!�����eF�Qi7tm6�u�*p���p��yRA�bw�I�s9��������ӗ��: !g��/��D�y,��5ivf��>2u�C�r9'����2��V�@����<��C6X��r�<�{���+�4Q�Φ������U�IA���?~� �jE'���]n�֝Wfӓ�@~��<1:��sw�g�#���#BޖUt�/rɇ�� A{`q�=�)��!*���N.8�L��5@�Fw���cW@22'�XzV�qn���G�s��j��=蓯��emW���z���b�f��ƯS������­��W�D�ݠO��!��#?4�Ml�˾����AW@�}��B��JCKK;����[�\9������dn͡Q��)�}H����%���2���ޕ�T��i9f'���;�]�ޒ�F�W*O������������R������sj�_�9�W�D����Y3i�S[Hؼ�f��Kijl?��t5���թ����*��t	'-1�\S�����	��ᒝ�{z�(AC�LS��W�gv\�M&@�|>9����~q����������fK��X��^�� ����{�=g��x}�r�׬��-G���kN-��:�a��xVJf�ϫ)���&@de��T�w�X���7Eu���� �*E�����v�f/Q' �%&��lJx��6�<����KY�3��Dk���~{�� s]��]�3�щ��8tp?$�4UG�X�����?�s�v��mrXg!,:g2��2�i;��$}������%�n����hkB�u]�J���Ȩ�M�*NV���%��'���#�3 �*]>���/%�.=��}��<�	��x��P_��q��V����z��(�%�����ƫ0UI^wѡ��r=�UiW�Ɛ�T�ОP�k��p���
�8��h���?�8lqn�ꦉ���ϫ2$�� �8l-� iM���no3��|Z�L��6?~�X�f��'�nmm�uh�A�U�/�C-�PF�=����v[�(�Ѭ��J>"v����!�ؠQ%��/�ʒ�̟|��@�<} �[�\��4 ��d�����;?�SO���`���
#ÀY֯�Ѓo���6]�m�����>aݓ��!���g=�D�:B8�o����2�G�����ɬ�26[#�C���Q])nY
�u�Q�A�EU?�|�^���Z�͖j���n��E��������ͣ���KKJ�e]F����/h�R�˅G#@R� �:���y��Qc}�jpH�xz=5��l�`�t�%&�Z�s�J�2�	�L r�i�e�g�k��Q���eg3����B��#�<w����U9�>�8�*�z$p�LJv�k� t��P�Z/�-=3R^�xk�w344Lm���O��~a�}q��CW}c���L�F>_�.��/Ƹ���u�+�(��i��{�[I\B�%�Ŗ&Hw���G�;4����X�]��
7�)���Y����xD�c_�0u��������M��j^e�/Ls;��t2B�raGo�p��d��I�D�Q��n긌�`6�Cm��3]�������y�8���s�,"��T�o��+� �h�Tݧ��o��!����x?K�0?:�����Sɤ��[��7�xv�͕Bo%f�G�T�%���^���'d����M��h���U��R@^�|������[-��HͯJ���zw;&��r��%m
s�2t,\<W�&G�J�g}�+���Ւl$��� �h����<�F��w�"J*����߾X�R�Q�@t��'V�xy��e�����~�=��V�JZ@�����oF��V�3>�H���ج�{��0���n��O/��i%�B����] ���z�@�l8Q���|�Y�"{��ng��}{�$�ʑe��L�:zy��V#�-����c���=��1��}/�Rnڤ<��$;��|f�%���t���������6�Rgo�ݍ�����s̰7��W��� 󜻜�_Mq����=A���⹥k�;vZ����s/et�}Sҫ��%��R�'Q~�Ԟ%~h��yX��,������*�i����z�mV��2؈0�ʰz�������H����O��i�Ҡ���HN�û^ L#k��k^U������Q��uڥD��h!�S��V���Р��&5�����j%�A'����Ǟ}����2�AI�$���)Og��&��筆��V�i���9�6.����tZ8agqD��)�VP�6�+fu
�1N޵^�F �gE��MT�Y���cys�6d.+��
�.I]�)�v��ڏWN�w^�h��N���1�.�ey�~b���F;�,�fB��Y���z����6s��L�hG�n-����Kd	>Jvt���T�k�̽�r��܀_b�6H0�k�S7��4�ߊ�⮰��߁��غ#5.����A��|Y�h�s��%<��腔���/��W��}ә^i�A
`�9�<_~��:�:?�V�a�k����Mj�dg�t���.�OK�\i4�'Wt�
/�==S��<�E)�oN/Ǵ@V=`��k^:+}���Σ;��ࣴ����M�}j2��	|��U�t����y��I�fF�_^�G��m�m�`�85]v6y���2wϱ�[�n)l<�e�c�5�y��f�4Nft��E��;#K�H�ާv���	P0udn��r��>&Q�z��+#���-G�jd���ٮ}z���Pߗ��Wl��q��|iW;��Զ�Ж���@��͂-���ã�u�Eσ �14�=|�q1F�	��?�O/O������}�Ǽ&u��4���_��v���b�u.��GVR�SAsz+e^���K�%
������+�;���(^�}���@+�"�0q�A��o�1�����|����F>��8�}'ǿw��������B�X�w����Fu�ܓg��%���}(^_*���r�Λ�8hI�V��Sk�[�NY��kM��%P=� �o� X9��^^
�<x��}4��l�@�(gb��ݥ��NU��"�B�䚋gyٓ��p�Z��L�z*hA��b.o�ԍΫ��[�B�-��U�a��~5򮉘�}�����>����q�j����վM�֮��ej}1��a0�Z�Ӄ軔��R��]d͵S��wn��ѓ,[~�8�](l�&�ɷ����P)y������C�nQ��D�t���+��d���>��#a��UmG��;i�^^3��)t::h���ڟV����3�� f��{�ӌf�7��R�1
�2�� G�I���s���Y�����;폆{U��@ͱIԙ5������ydh��fV�)�򺰓�V,�49]]!�_�Fɂ�
���Iӧ�߰�rd t���߻�3D)�Ӌ�2I4�z,�U?|�e?��:���	M�����{����O�^��<�j}fB�Sh�sG�Y5��K���hÿ��/��e6��e���	n�z�g<ɺ�
ʴ�|ޡ^hT��¼Ϻ^fgL@F��2Ԓﻏ3}j�iP�`,jT����>���WzAsV��J2�A�`�`4���K5��W쑉������$���,bI.7�Yr���h���w���(~S[���G����3��8������yH�d'�*�	i3�>�X����p2���!ڮ�m����~ֶ}���j�Bc�-ֹl��ΧZ���4�E��h�����l��������t��)�+Ҫ3i�hL��+Df�.zHS$�{][�C�*~�}��t���@�kZ������j�|;g�����E=y��v�[�`�eC}]c��ӽ���"=��	S����u��^�Ԉ�-x�r���]dh��R���� 9��ހW���<��S�.Ѯn��><�ߧi�\�Bm���^W��ɤ���?��<R �M�U�-�������e��{�/5ʔh­�pOj�\������_�o�5>!΍�D��@9�Ǟ�]i%��N�~�5`�ϸ6�5�pÂd��"Z{Ahg�:��=���	s�ó�"��>����o���?�ۻ��-�׫�x�ƴa�#��R��=X ],�R7<��[����u�L��Z�L�N��X�K���Ǡr8O��i��g���>��Pu��:<��䂃c�	��I)�N���.����u�g����ǣ���\��x�Z�J�	�����|��n���ėvO|�]��ﹺ��<�vЪ�?�Ζ�t��)ߧ2k>]�������E�Q&+�

�u�!!�I����++֝ɢz�u���%��Ӳ��.M]�x4�sEţ�IA~~��������)+Ƚ׼�����)�7���2i�,R�A��4�)@݊A*�%L:؎Z-��5R'��JL� �	r���3:�s�E�<'*T!�Zظ��,�]�f��Ɠ����C�f3=���el�ڕ�
��|���ֽ^�эN�'Ĵ�OV9^���]���X#���! f^s�/���+]m-ɜN\%M!�� w��Z��`�!G�S�]�u�����o���b�_�o������s[hSdB����z??6�ð%�I�� aZ��?Ny��
�Z,���!nп��A���jJ�-��S��3�J?�����S8O�c�D���+ǟ)�8�=ݝzO0�e�yaр�t �@��n�/��{k��;|rY�������KG��pSIf P��t-Mu�ɇ�&ߏp�L���	r����˛l|#��ӫ���6�.+՚�����ǫSo�Go�&߇	Kj��ưw98�%�b=rr���{�:�ϻ�\��k���Zt���Dӊt8�RU�#b ����hI�Q�!&��Pc����L��g�є�-��RX�4�����Ԯ�x`� ��F��oQ���$���^�u^+�t}�W�`c\~t���m\~f�ӛ˴�l����u�	Tiu{o����#G�|cAZS~��A�I|��D�mX�7�xc4naw5l��N���y�g�yIp���ܜ��br�A��d�T�Mګ�IӞ�O�0æv"�;���u�{�����}���#�������"H���w�\��[�x�@�rF�U�WW��v�&{�)�O����<��-RRR���9o,�A���4������H'��xz�r�\��&��Y>���-)�j��/.�G3��]1ZV���B��J�.֟!uc�\����'�V�ar��B~ʖ������2=��B����E��~�<��w4��u��ݝVHIZ�ÿ�8��<���ewz-&�Yz����n׶��җ�4�j1��iU�-��y���ƒ�أ�^I�sEF�"�ܺ�F�o0gւA������}Ɲ�9�G��+��"t��w�SRZp@K<<&(�~��o҇	]S�)P�Ë�:��B1��m�����Q�[A��ot�~���1���k�X��Li	-k�r\����r.��%�Y�Vw�����7E������^9B�NB����"/��H�������C{��'
�)��$��c����zޣ����M�k�& �ħ7>��>ݖ����n�F�8�T����v_���w��m)�Mo�`��zH�$��6�;�
|xc�������<���DM�S�_�����CE�UTx|��#�L�C]�-..�����@����-������g6�I�",��(�������5 ��R�ϲ�qdt9��8u�%5��'&9��ܟk[����E��
��[C��R�i[DT��.(�Ͱ!��?�,:�S˺/]VsW��z����B�c�hzHO�uM�0)��dH�E��N���R�
��a�ChU��^�n�y�C�/u�;𺹵7.��ac{��#�j���P�tk��1�\^��]��w!�rJ{Wi��9������cČ�F�`�(�;ٟ��Bw
��� ��γ�Qt�r �	�\[��:~���%=�d����kY'�|v�_���kZ.$d/�Ƕ���7/.��d	�nq;�
콺}5o�-a��=�K��N<������Pw3)�«���ܠw��v�ߙ�P��S(���C�t�ٓ���q�3��dٜw���{u���A�(
6��5D���_d7f�����L����j��m٨���/N����ki��_����J�dկb��9�{������+BC1���b�슓���î����I&�{�N��G..�*T����v6��N�n��zO�v5H��c�BOb�7�����c��fJ�5"��F��1���\F�u�5�?�I�\݋�n�@Hy���Y����ޟ}�vVh!��%/'%~Ud�r�"�U�݃/I��XR� ���0T�^s��7���ϳ��1��Z�[d���֖���C������2�^&BTӽ7��燁-<pGXț��(Ee�$G�j�����I����Rh���i�W��s��k&��f:l7{/�s���g)�Uȧ���Ǟ���u[DA�s5���3��Ι32���8�q��bF��d���1�M^F���n�[���e�tN8���p�^NAauc3Q)k�r�၄�;�T�O��й��7�XXX��W�jϘo��I��E�&@�5G�<]Kw�ҮlR���F�tO��W���3�g�`�R���h�]o�,F<L�r*^�ՙ.����_2��r��W]3�Kb�����C�=�s��,�������1܁&<��5)m��'�OG#�63??Ua'�$��2�khs�?�R�<@km�`z5=��܂����ԛd�Ws�P�Q��\���CϦ{�=\O�&�E�STQ�(��J.����,�2�%���KCX2����c�!��0��/������v>F9�AX���\���7�덎����kW>�iem���
��JˠRr]�>L��� 
Q�f��ٲB]^�9Y�@�*�N;�+
:��eF���̙y��	�W)�'�r� ��$����䛓}�(�r,�7��q�+�3~T"_�zg�!���un9�J|�> 6�����@���gc0��/��~z���Qd,��xB7#bn_��Q��w�&9a���D��`��y��36�#��Jbm�w�ne8^��¾��p9�\Q�A�,�����8��(W�_����#�P�І�|� cF,У6����Q�_v>v�X��=8r��YX	{�3q�/��iX	����1���f��q%{� ��J����+E�{�&�����=�A��OC����T�50
��7�*&��ԯ���g�y���٩h&*�>z
��fv���)�h�"�Y�Ol���������0-r��/n��ʬ��j�����F�!�I#s]ޢ�:#6�7��+���\��r�N[�������P祹�|���߼A�~a�L_ �au�0��v���������燛O���s�a�U�t��*��aNA�E�dH�%�Kn��t�T��J���w��2���a}��ǯѸ�n���}����d@��>G]�y�b':W׽�EF�z�7~pn��7���0����4,�6;�8f���7���x��($�1-G�7�#��,Sl���R��1�+�E}���� ���#�(K��}SM�U�Q��JVr�;��6��w*�m�����O�ى-����x]���.�@�������k��?���p���%[��ն)$%!*0�7�M�u�2�i�8*W.��A�wh=���)����r�sL�֟�x����¿(��X=19�lJ:�
�T�����b*C'�
�I�''E�_���n2���8t��o��2����D��8]}�]Pߢz�;&�����}����+�|�JO����*�"f���ǍV-�b\�IWq��,?���(�DJc���/�����\\�i������H<<��s]G⥥藝:���l���= G�
ʟ����SF	���2R�{���_juu!_k��d�p�u�qs���D�V�.ZC� cZYY%=��_(����>t�\ۍ���><���X���.�#gCũn��+�V�..��cP� ��=���ڈ�� ����l��:���*���D�TCj�\���jfϪ�'�55O�C'1�8m}Vjt�o5^ߪ.B7��j���ӣ���gV9�Y�׍r��D�W?���\�bM�/�9�mLP}?�V��ЦwQ[��=�c���j���oHm��tu�ƽ��z��0����H^�/�u�%����`~��)�[>]�����m���%�$��a.9��y����aB>'�ͱj#T�W0撣 r�2�2-b"�2d�+����yY<�^�UG�#M�v�j}_�۶H��:G�l���(��!�����ν����%��m�z�A>��9
�x���|:�Aަ�u���K!�k�ulst#��[�h����(�t�_�NG.W�j!���ܔ�]|O)N����+K���zh�������a	I���7����&L혵�\��]-�2�F*s�G<.+
0_��u'��Þ��8��|��d��Lz���z�w�.`��}�:3SZp���>�����|Gb��g����g�X���y�F�������S�d}_p�3�P�e�R��K���9��jR�ӹִ� ��5��@��^�C[���v��
]����d%���S�)���MQ�'�6�1 �j��t_L�[�^s}m��U�]�Z�}klk��E�Wn����l�_l�0e޲#5�AH�¦�`O-Ze�?*�m`�8��f��r�(י�4i�7���8����Ѭ��~{��(�.�x�5���Ȃh��Ygl�Z�P*b��&�M��y��u��i�?�����(?%�Js�j)^[�"ٷ<jתޒ��|�`s��N��O��N]�w~���ϙ��U��G�u���s�e�l0�ɡe�5lq��T�f��/�
�*ce5�D�L��H�+:���n09T�x#�t�֎�}od�����Lp ~ɺ�.�:g�{�ǭ����M�Bg���[����.�.��K�L��L���QV0�I��p�{���q�d���ǫU k�o�d`��M�c��_���d	d��2��L��R�\<�	�֘}i��)�������cc��M@7/�l��w��B�]�_��"H6(�C&���2!�����Ӫ��wcm����5m8��$�+x�,q�qȈ:�b�~ �]-t�:��ā��e�o�L�TET9#K�(���a��ᾄg�M]ljr�\��4nɕni�j"�~�5�%ơ_\��{Ha-��q�uE���TF��PG�X#Cp��`c$�<�g �}:f:o��%I�<�kLԒ�q_%i�Hʙ�c�׳��������r�k9�0���P�2S�,���ox/Ӗ��*ч�NTnڊ���/DZ��7�p'��T��v�ctU�ba����2G7�{;=OɝWЊeeeU�h~�s0]=�=�C!�_W�e�i��t�ϩc�ߌ�x]F�wJ�m>��յ*?��Tf��F<0qn�q���Qi�Kz~��a�<e�����j1��i�k�#�b�at�4�@��� ��vD�t��OT=K���Z�^KF�`l�Ǝ��e�1T�	��Y���n��*���9�L,bY���ڮ���qiJ������M�{�H������c~-�k������1(N�X�X�<V�(�V�w��<L��a��_�E��]z}$�Z���H8ӊ'��i<��M����"��OG�����׆�Lɺ���[�o�Ą�F��{����/���cߌ�J�e���6�l���6j9�ft(k[�N����;�W������v3���9�9�TPN�32T�������
)sZV=ZV�)ֵ	�'� �Pm�x��e�s�GJFV�����T>��U|]CG�C׵+�Bď�lGKH&�����Zw�h[DR~������: Z�&)N�_�?h	Z��G�R@��Y�P==Y���ʲ�q�<co�����`#�o�{�pڬoC�Q3��j��?�Qu��{d�;��.E��v٢����M��敳Sq��u}!!�p�~}�-O���pg#����u� Jc���NRV#��$����$����0�R`PP�{r��g�]FLݎ�p�O
e��X�ؼ��Ҥ�A#�rj��h@�PC؛,W�{]kʚ�s������<���-�K��+;�|]���uJ�G;J�1a`K>�d��D0fE;]c[���sl�j�?������]o,�?SG�����e�q�j,��N�Sv�%��Qz�'��c����@(���V ��vV�b�(��n#@|�b6Y��BU�����N���,E	B���2��!cJީ��q����L�=�`#C�B�W�
�S�9s�����=0�o4�w�q��/���1�p ��&�
�3��F�����+/������=v�Ç��JZ8��J���Vњ��	r0��ki��)s�G�i�jFmГ��=}���j�߻��ގ(�P��-nt���ML����X~���Η���9�o�y��(݌/�����Fޔ*.�M���id$ƣ�;�7��E2̻UȤ^}>]hp`O���)���r�,.~�'���)����1M;�dW˷��^���*+)ss��u��m�q�؆��	����[zy6��8�$�W�L(e]4�;��j��*Q���Tʄ�I��gD�l����SV�����JlQ��;Z��la���.��Կ�#���kd;�.�f������w�<ݪ.ӄ1e�!�m΅\��hP��n��?lV��N�3�	�,V���eS�V�݋t"�|�/�{�u8������
RX@!�oB�%��m�]����&5��C�C�e�i<H���?	�~2����ޝ1�X�H{,߱B�񄅕0��դ�۝[{�5W�?�[*=�7K*��5z5�n���$�!@���?;����}N���1�PO�4XT�)�a��>���p�u_�����\�������ʀ�2j�H�����;I�N����o!,..�Z�]�T�2�*���!:��O��R���5p:h�17��.o�J`������~�P�����~�]+�^l����3�&��fAF,�Zf8���y)�+j-��07���w�'������x��8�]�*���|-�U�+VF	�'w®P^�r���SE.;�fa�F����1��$3�L~̨bi��$��1{�C��\�P�)g�o��$�	��;
�����_Ll���&y���Έ~1�Z|q����+'K~�����ļ�/�E�i�����yV͆G��@�p�p�����~�w�W�,�i�k�<�amiye����m�������r���%�`sH���n@*#�p�r<ot�T$���ޙ$�e/��D���:�E���� �F��������怸!�ͦ�U�f2|K�o����	{����o��_Jk��_�*�MTs��z�l���R  �5�	9���4�I��YG�S�zv�t���b���G�qG��`A��  v����2�|;����ZA�PC#ê?��0cQ�g���-X᪄��}v�b'զ�_�-���9��8��N��0�k�^�&�.k��bf��]�k"c��Rk100�t|���)x����BG\ګ�S�'�onQ��q5
��(T�{4^{�?�zĞ�d3��O-�V(��*TL̄55=���-}����J-*R�{40��7�de;��z�tSt!�u����s����8!����Y)C�Y�3-t
s �7��C�G",,,;�2�Z�4c6 TY�,�9>: �Mv�w�5��˼�`��Ff�]ܨR����J���?
i�KQv���7�}������ ]f�LI0�v��H���2Tr��;�KM����W\eЫ�^�+[Ŏ;k��Y6�}\\ί��#�`�&>Js�ظz%ؤwu�ȶB3�e&�ȱS`;w�+ۉ�E�4z����.h|;�g}� ���Q�`�?�o�^^�u��x%�{����5�8nP2���*Z-'r�+)o�=�l������r�<��u/�<L6'�S-U��*� �V�Ooٔu�tHQ����rq8~0��D��dt�-\�W; �ՔPf��=�2]��ܻ��Ԧ�vj�<+�����wÙ^���w.��l��p�6W���q9�,����7��w�C֌7g���`���u�ǵ�\�EJt���L a����l����~Í��a��㸙DǮ�2ڄ\;�����p�s;����^�çx����t��(��\گT��D����F��#,�ҥs���o7@5'��[�Ė�S�f��������Fr����fL���Gg�L�+U	;��۫�]�2���f������(Ӄ���Zܱn�e8����� ��^�2�lI�?sxt������O�N�H���o}����2��%����!M�����	@ Ļ#:��7�TTB���<�/>=��7�� ds�z],�Z��H����
�M\f�;���k��Xw��u�G��B�ID�T�@:~?�aAis�����555�	�T}�=���BP�TA�#p���������۾��om�:p�?U(;�����7�m�,��N#Ϋ������D=�Y4�՗� �щ���~>Zo���ݡ3j�"��"�r�*���+��Q�_��hF��2E���b������;�Ե�7��H>�b��r*���b�v~ `������*�S#Z�ݦ���jYJ�f1KtO��v�e�ݘ�����(;����� �,�:Tci�u�pC���q@tCjIP=P��ˁ�Q�7`++yP'�P������)��gN�/���sf��xm��'٩Rm�!��$�*����|�{,���y��Z���F�а  ��U7�Z
t��&s�]��ew�{}ď�E�;�tk܊���٥����O�O���u�EPۙ�/�w�F?�j�U�rn^A__����Ol�3�ȴy��z��b)iX�J��b�Ω2���%9H����x?�`�<Z錻��X�~��Ғ��V̫*�K/����b�*Co?V��#00��X#�=3�A	`g�_Nw��6_~����.�ù��[!�Y�z����
���ڙ�X`�VTޫń$��a���"��c�x��OM9��w��q9�Y�$N�(¨�9��PW��� ����`A��J���������sϞ��3�t�
m�܊	mmmό��*K�1�[����פ>�0&���09eP���m�(��*ܰ�޸�I䐞�  �s;��缁Э}q��:,+���K7�*�����h*�10f���)�HP����=�ߥ����D,��w�q͗eA������3MV(���O����A��ul�� T�6jMv���7&|ƛZԣ����$^\ QŅS=�!/���8m9��}�F�bE��6d�ћB�����7W�?�}Y?�,7=t�\��N�տ�u�v"��U ��Z��8hÄmh����ҋO�fy^H��> ��*.�_F=z�F���hΣ�o�iJ���C��	O��A�1�6���A�~F�`C�B��3=n{'�2P���c'��D�^�9	A�Ȩ,�S�0�&Bf��x��\�S��U���F�qBI�O��{�>�9��~�s��^���Fը��N�V�6�j��[������|Xږ']0�n�'�'���}Pf�s˓�8=n<V.s���lV���JvY��j>�	��ap����{⋉�s�MA7����E0�na�?[��.�K�?,��5w�|D-���ޅ/����?M�P�@(��-�P�ԓ�<����`��C^�?�ÐWv�t�_��3q"$xܮ��`v3��S�����/88��̞�(�D��Q�s�; 4<�,�+lU��M.!aԶԀ�Z�&`�"z��]1��+���ʸ�j�`jݓ��}_��XP�IvI��M'aė����q �t{cJ�l�����Z���`�Ea��Y2<s��,�8��l�i�����C��
�onvg[C��tv�#1�J�������k��g�N�_k����Y��+A�<Ų`��LX(@��W��9��-��Om�,�����)�ֶ��	P���Ls��Ao�­����~���u��HТ1�����T�`��,���]��0���_�M`U�7C�#"�;_{�����,�K`��}Ϙ��9�� 4��r�q���AzǦ���L�Q��ɱ�����k_�Q!�	�	�r߉��zՅ<Q�ܚ���CL�k��"R�V-���(� ��rɃ�A�lw
�Ͼm(���i�����_q��:Ӫ�|��b�3�]i!]=0~^�*�U
�%a�-��a�����_F;�/\tŁ@�y4z'�.��`�O?�/�z(+�Tُ�gB��� ����i�QK��0 ���0�<��n��{Ҕ(�pWӜi��u�ӋEEb(��˪Y�igH���
��W����õ� 櫌�*��̨O�FF�>�����>�$����0���wi8 l��wJ*!Wӯ�v� 	���-ٌo�y��{��c���_�_�ϫF���ge�V�!�FW|'�\X��a�49���X�,Jj�b���U�����6+��	�K�h�sO����# �Oc��^(o4�m�9CM�Lb:7��}��/�Z��Q7�0Է��Oٽ���zr��uv��֡�H懖F:7��_H��U��3*���NVڤ�t�%����8|%>�ĵ}'�o4����h��0Ƨs�«���E]�S(.�G/���ffJ+���.B/�S�ݨ#?1�����!��*]h�;0���.���'m�J�G�� m�u���{�X�N`5�q�t�ʵ�SŧT����~7 �%����q҆&���,�P�O7:ފ��hߺϧ�xܞ�^�eD�����Ec�<+k?ou�����s-;�|�m��j,��(�h�{��-m�W ��E�-#J�r�2� T-�ۼ�����6a�s�er�s�x6���9B��d>uf��m�]�����!��E[�ןK��N�,R����e	���(p��<w8�����R甪�[�K�qn�'�U_-�$ɨ�� A%Sh3�d�z�x�%�L-Cw)EEE9�/�����fpBkT���ڛ�r�*� G=��I�������λb��K#���9�4��r�w�α���Ԕ���u���=��Y���[uZ�P��H�6Wh���&`,�'U���Ƴ�S@1c~���g�M�"B�@_�swZ������l��i��k�?՛�~f%��^��f0��;��6�o����ec_��j&���z~[<����{�n����H(�w����A8��tӽ�ζ�<�M���S8Fݦ�%���Y����o-c�b�)�=
���X�Dn�g'�Q�e'&��n/� �i n6���y�ZXO�Ԓ�\�����V]�WUW��N�74%�\aK�pa�9&�LnΆ��f���!v<��Z���t��sN��(�ܟ2��p@�!v^��"�~�Bh9={��z�YW�1��?��j�***
o���h�۹�\�=@}�^+�t��i������&�O��N_[˞�A�Gb�R��Ƅ�t���>?��)�^Ku>��r�\�ƭf}���ْ������{����=��-���e���e3+�2q��T����F�Gϡ~[0B�Pc�E��/�?;�	�w�A-���84�� �6�� *��_�*��H8����L�����T��Ѿ%�Q�S�J����Jfje+y�j�3�D>AY�k^��^AGJ,�E�tj�Ʃ�^�m�9#5	G�"��Ѳm�����%��;ʛ�t��XJ=��#i���n��nI*�\�Fؾ}u�4�	��Ν* N�h���v�	�Z�-�)j�+^m'<�|I�I���ٓW�%ꖘ����B�*��Y� ���	���=��'��f��Q�S�{����X�u�ow�x��M�0F|�F�,DWh��U��ͅ�+ࣀJ��{ ���Pp�U�G�O:����a|�8�ҭ������[��螧�Z\�<�_W�1�s,_Y����gl�qX�
jt��$��<�`��c��	����"W�? �+Q*���>�ܿt����.� ��J�M*�����P:`ɶ�*�$'^bM��)������Ri�ؕ�?���8�J�#Ϯ�d��A�a��e)bO��S��><�ߧ�2�̳�
�*���L�ʱ'T�W��u��������X=��7���S����?��	��y��ҫ�?��<���W))q���!Kٳ�,%$!{���:&*��d��}���B�wfƖ}���{�fL���|�S�xm�u��<��:׹*m� �����z��y[�9�5�~Ͼ��ͷ�gJS��v�dzx��Y���P�dL�E �a�¸����ܵ�[M��\���{�?�).�Rv��2�'r�qS�خDI �w֦�{*�p�>�\+T\�I����zM���N�|s.�7%I���8�S?�^�x^Vn�D��;�٦їG�F1ʭ��}d��I��e2�-������V���8p���>{Tn�5x���|�e������A�r%hPKeuq8�E.�$�d�c��z+��`����������~��)��Zf 0@��~����g0Ri�|O�����'��B�S)�I�?���%c�iK`���dW�(���N��� �G>���O��t�ȇ��w��׫e?�C2��<�6H��*�ѣi�Q�Y��]��C"J����
�q�	3�|����p�������'�ҿ��`�E-��w�D��8g���D�������95�������Y�%x,*N��cs�-\F��/��N �!��>G�QDщu@�H��ο"c�Z�2���-�w�A�T���z�I];�!,�� y"E	��H��;X���-O�F�R?$���P�;����!b�e�_��1��6*>�{�S���)���eP�y�М�~O�0S��Z����FF����[�u�@��јj�&R��r���
9���h<��/S)�	yL)0 �[U�]�#`ce�}�`�!����S�@�3G���4|5��5�%R0���!�6�<n#ȑ]l�y�����E-��㎳c� �+>Cɘs^��1�����Z��!?H�o3*����h��N�|��Q^����V����{���/t��C�|�n��Tk�_Q�v�DH�1�ϗNF�uG��1H�?qk��H��mKL��(K�Hs@A�`˹j�>-+g �[n�~��:��9�N��܆��tui�f��a�l﹪��� TG�_����jPCCK��zb�͌Ư^GHV�{OU�ͳ��\ܡ� � �EC�M��2e�s,�{!�ʽ2��#�I�d�ܻ�'�0vM�%�ybٌ�z��A{����^t�ko<�"^?�.1�Tܶ����%9���m�[�`dWy^N#/�6��}y5�ڃL����t�ǥG7�sj�\��������d��I�������ߌ���YLRo}���HZ8dejy���[�&_8�r�s�q{c��,�x7�H/H�f�l��YN��2�[\K�����D�>���{�bL�}b����|ڛ������c2ɍ�]��x�9$CFU8�% c1 <����J����+,T��g?N߷�Y����m-�Rp�v[fS�����tQ���P��j�Uj�x"_2�t�&��/TT`"�ED�:�� �8vX����.���ԽգC�jU�00���ěx#DA]ֺ:_�`��yг,p~]*�1SI�U��e7Ojݢ���~7���۞ۨ���ȑ�*.�lS�=����?MT�&��a��<�{2|v�R�#'�;~��9���G�X�t-I����[F��l�p�o�D0X��Jިy�$�y<���)aH�R_��?J2�]��X>�]�D>�����p�@����wߜY`g�}���"0��A.�Nު��g��dr�V)�SƼ�O�lO���I�.�FP<�`τӳ��)��R���l?%a�OZ�*Ȃ��U�K��pi
�b����n��gK�-��V�=�P���\�|4�`.��H��y�s�0P����/����p��M���w�\��NI2��4U�5���&���
���L�?fљ�̘V��k)��y����������*��k��A����]͈2G(���G�w�� "<��,#�DQ�(��I�d]v��2#Z�8���B��`�Ȫ��v0��g#�du�|�uբ�����/�CI�`Y�̸`������0��Z��IC��o��5�em���7Xu��3�.�>�̴_����־/&?<���,��f�� _�P~��1� ]/$�Tx��k_U[^�B�dM�<R�Ol������i�t���o���n,X=����.'��r�6�\��Ϣ<�W��S�I�su�G44�b_�\}�S�1&=
��W�|���)�?A|�����LQ��4��H���6L���:���NO7�=����!�JGS3��P��RՔ�|�j&K��7?/ƥ{H��&����뙙b����7�S���~.V(�}�o��~f���:GeI��g��~5����.�J�r'�D�n�N_��ot�����h�ތ��@mXQD��p�?��`��\�[�I��#�:TZ���=L�t�+BF�oTg(��Ar8�V�雔�{NwAW~�gƧ4���ƽO`e����zN�K�f�w�� +�N��34��BQ;o��<�����?��i������t�o}`���įBbT��;�����۶ؤ�[��A���1�
L]1|��U{�Ճ�q��54d��%]��"��zD-���o�(�]���#l)vg�\��k�� \c�����?�8ն�܅�wa����|�gxNU�%���"��} f�9ts�?��c{q�w���LpS	�{!]1�ʋP������!v��o���#���P�1&']�F넼���}ܧ��W˳,d �6���ot�zjf��^_�`�e�uzG��f4�Mu���|o�]�R��c�=q��P:��&�����tA�%%��dvR���"���ZE�&4 RYWR��K�ϋR����������]��a�X��U�s~d
��,>a��:z?~���=~��N�r��\��Jc`z������m4 ��n����>��5Q�α:��1Ddff�ė�ݖ��x*�{�$5�&��f\�}��1rLx�Y�U�4���7�͙�%����) ���Pã��"	����+]7ǳ�����hW��G>͹�\L�ώHz�"Ƅ��m�(���6��3I���W\<�<R�5l���"��?^�MaF�w���&��b�0���2�����z��0i�v�����D+3��U��מ~��}�����Mɚ@Q@]|csۍ�<�0�<�����+�P�ڵ����R��
��Q��l�v���n�6×��3>O�;:�4������������G~t�_�\Ԋ+_��Y�G��0��So��_s����k�ڗ�ڥ	���?��.�t�S#�ZunX�C�AP_ڏ�h3,��J�Jk�{~\5.���`s�K��$��g�i�`�\9c��Kٕ��u��؀��8��N�xtj�J����P�eGW]n%ڡ�~F���`ک�sT\Co�o$�!fi;tJ���I�W����k��è�\��]�#n��>��O���!+���� XM3��)`���O��������q��;&��?hν�w0Nj��L��GCtc����r��֙;R������Q��T�R�9� �L�	Q��'�)�B���t.J"��|;�hI0�MC0�����Y�"�S��`\��)�Mv�b�����D��Uw��NM#<�wtP�����m~�ff�p�]Sҗ*�Ջk-7Y�v�0>{��1qgE��
�;U�xZ7�d��D6�m��n�%~��j�� �,�ύ��g�7F���,�X�8͞ްnnm�H�Kz��� �y@|ۤqW�0�T�aL��c�غzX�knq�d���i�]|�$N�I�*�}�m@+q>�xo��E!|��AR#a���|�p�Ϡ�[m����<�vA7��ڴ��n�������E(�Q���䧞���S��/�VUT�1�x`y�R�ɿ�� e�|�g��6�Ω�R�D�^�I�!M<������8aM�m���r,�g�u��'�]����rO�Q��^���z!��@
:6p��?J���Xs�r��%f�|ۆm���M��i��3e*��{�S��c#����uf����ϡ�����X#u5�XX�rU]+ ��� �[�`Ø���q�9҉���腚��>xÁ}�*�����4t��ι��~V6�5��B^b����2���/� Z�� ������J�J6�'�������v�����YRNIϧ����w��c ?Op�n�_()�f����B��
�fYm]vU0lm�d�Y�R�ɑ�Wԡ���>iMP0�|ҽ�j�h�k5�ayd�| ��o��1D�^��TH�b�Y�{��p���
kB�}N��$�<���ҫ��i��E��"�?)�Pňz��
m���y��^:���|��7�1Wf�kjH���휯S3xy�m��R_y-�o�
cu�������0��F����AMi�H��oI  a���1��uPW�����w�9�a�L�����Hg�n�uO#/�PZ95�����]X:���N��(�<'׵�%E/�#�
¢@xns�������_ �ě��Ȫ�e�K�
H�z`�K�`D�/�DO�jY��+o )�����oީKJ�v�9�8��\�ߌΎ���<s���&��K�]���\��pR��>r�6>����ⳬ0�ȵ��w�H�,ٮ g=k7�������*�z[�u'�P�'�Qx��o[lH5Q���2J�p�e��+99%A��{� �h�=�@���U/ �دcP�V()8>ů�����Er�������!ʛ��ĝK�<�(��j�Yu~���x4O�2�E�mZ�ښ{(�����T�TX!��9�K��,-�k��P�JNo���u�>&�d���x�뻪��έKm�e-�B�q.�Qsz�J�l���r����Y��H
<]�I|d+wv[D�O�T���x[�i�p��2�J2��Yo��_"�<��ȏ>������y܂��l�D4xk��m1�W�O��kh��)&�����2�^@��Hd�e�<����WF%��2������-P&b��"K�{{ٌ=l���1*iR.1-+�C��?8H6����7�y��]�ͯ	�7P5x�E���Č�\�n�[.�<�T�?ɵK{��9r(5N�d|A	;���Cyvv$�����\�^F������#���`����O����,u��օ*o�
¯v�9$R�������F`�.mK��`���q~O�x���6Tқ��ΝP<�go�؏oӐ`�f�9�я�x�
o�<�D�=�z����Ȳ,VIʔx�$9Fo�N44�;ǺZR��U�&�GV��-D����e/�1��ڷ>���=�*`z}r�]�`A}���Y(�ܸy�����6��5@z���cQ��V[yw#�:����,��Ťܤ��J����Wl
�:�?�o����Z�mp�����<�އ�O�������'�]d�s2��N�=x_�'I* !�#M@��+���L*���=���f1��������Z�ؚ�����3�LQ���TO\ސ{<F0(,r�����8Q�^�2��1H�ݘ�/+{BB�~�r/؎<P������9~�m�;%��8-���Xo�Œ�����T'��m]�Q��,��T��?s�;��B�\��X�l�x��خ������ai����~���<w�(� y!��(11��$\H�f��Ό1�!i5'�S�c��U�W����n�sQ�æ�r�Xէ�;̰���7'��<v��"@���j������x'��_.��iD	# :����|��F��Ξ(�H�o����<���%8���r��V�6��4D�h��'u��nB�
�m�S�8���ˣ�.ߐ�,���wL>e��Õ2�𐏊�7��9��O�`C�n�W�)H>!�����YR��!��q���
�j_���AD*�Q� �+%���
��������lzRV���^QV1�m9&��?+s����e��g�p��mٽq� �3R�8!N�f�"Og��g�����ܬ��3��@�=�8������-�����:`Xǂkο�1��.�{���YA7��I�ڪz\r�n~5�sjn���''����A��s����N'�}�C! mp��������scFv*ꌏ�&(S�y�D�0�5�/���$G�?>\>%���Co�E�,�X�ɩ�yݔI,�U�� ��@������a(�ҥ�*�9�x�M
W1%���� �"�9�y������W���q�FVC ��	���,֖z�e���'1�6{����i��0��	��=I��e���R覇��ĩ*N����a��L������d�%p���0�G&�R[�6�S�a�:�o��8tjEx�� _.0�[��^���㸬�ԕg}��vk����y����03��xФx��`���䇤:�����.��:X�7���|�H�W��R���%C��_]�۪x23"�h�c��\�}z}y�5"����U��ِ�Io�7�	9uk�c�m�;�7��i9���t�ʹ�=�0t�|YVn��xO�~+e����`�	��Mgp�B���vԳmn�����t�����9cWdL��q%?�H;Y���h�O����w�&��;�E�|��)pma�@e��ue��+h�)��X�]P����&��k�����[�=�����[<��}����j5H��ǬR��s_Q�^��_z.;d!bv�.	��ݵ�Н�E���>$�|����$��NZ=��+���������ʪ�8�C����4�l���W��]��/�+�e�3%��4�b��E	�%e��/שO�����~n�����# 476m��<�i|�Ccݞd'ӏ7��6߇uLXF�'y�&��zui���x������u��w��{W��G��Ȧ�0�@��5Uȉ��rx��$c�}|��i0}�Ÿ	�!d�`�*�m����_zj�֘Y}�v%����~���"~T� +�!R2�]ǅ4J�Qm�M��m$������u��q�4V4$�:����V��?oo�?��C�mWFʕ����&��˾�%��U��� U�6�����SK��l}A3�t���X�$�f�D"����Leׂ�7���W]���G��׸G_���	�.3�-`1ԥ�\��b�#�1S��8��_�pK}���g�{�A�(��ufc���髌}C�>u5���0�)E���2��P�\a>d��_�b	D ��*�~�d����{��D�戳9���d���\�#�p�[_�;(@Kq�����D����v�����ނ��nxQ��ï�i=9�E���ag���Qrn��z��^�_l��B����y|����f�K�7�||�&I�yp%آ���9P�h�k��ܗ�ϻ�]��B{?^^�
�-R'���#�pc�=a���C�b���s5י#��W�Z�+�j0���)�zv�Լ��ńa4E�\��(l�(\O�L���KLKcj���S�"�����l����g7�t�-&�X�~��[J�@Z��~�[a�����cy8���7�{1�<�ޠU�Ǫ_q�S-Y����b��%��k0��j�}Y�q����ϥ)���!� ��`�s��^�<}�0ܽY���j׹s+%��.�g��~l�)��S}��Z��)���{�ٛ�G�>	�'=�Y���=z�V)�o�e��>KW���݅��7���䈹�q�Y�]������~����`�u_�H��'M5��],�^b�Uv~�Zf>�T=�N�	����o�m�_u��b [v<�ׇ|O6����(?�ߍ�)]�X�&O�9CQ���܋{Y:���>>����&��f�qW�1~Y���}�Ef�D�8=]�)�߫ƾ`�X���ɽ�c���������Q�Xb����.�_�#N�؟
���)��C:�r?�r뻶�g�bQ!,��XY���F�������z=�}�
��3��"�X�ɫg��u�*��O�m}t�c�Ү�/��ɬdC\�#���)}�5��!���{9�ح��:�G��`$�PҸk����7c/q��|��; P'�,�����μ=��%�h���5u�Y��Dwۯ��P��T��`��s�
�:[F��E����H'� n��W@"m�,��[�_'5�FFr��A۽TZ����w�����[�2�jޟ����.T�lf|���KϚ�bj�B�W3f8:d��k���!Z�w��6�
W�D�c>~��
��q[Ȍ�KM��,��pP�P�����8#R<nv�/*�ƙ?����[���A�av;������,Ά����iD?�'�������L�h�r�?�Ц��eD2�䯹�m���*�7�����d�'�P�೸�4�L<���:�E���g<��m�4�!:�a�
�6l<=?�U�y�v���G��R~~����j�s(..ch�ڳ��qC;�X���ܼ���8Y���|��\�LQ\�ǥ�N�����~�`?f��~xE����_(�ğ4-�\��)�·�˔Aa���ՌTg�L*�)�^�=�,�.�xE�p��E���� t�����w��������J�����v��YU�x��)�ػXw�a�1*��2�{`����vG�S�L	%������Έ����'�*r�Ԩ��.����x�����E�2�b���1���]���QY��;$ ���QHG#��S�8��E������\́]��V��a嬺���gJO"�y�Q��b���Z����$D� W�ʼQ9�U�"Zd:=-���UB��`��j�O"��e537noez���ڒ�d}͇���k�\'~O������f�fg��k��ܲ����;l��<�eb�7��D����oR8Z)�\�י_����;T����c�DE���k��)���M�����ru���BCR�[.�3��ڵ(��j�5x	��C�{������պDZ��t����Nv?��ħ���O(^K����������wd��9?��C\����F�~곫��b��Q���}�ڕWtœ�]7:�+lMR&�y��[Տ?���YQ�&��76Z�.e����_:�;YVL{l�]�1L�Q�R8��i�u�EY��m5�ؼK�O":ē��$?o��x��#K��z�^���7@l-Ok�<3��i�%���_H��3�'ϧߪ�u�_Po���ێ]��y��I�����\YN��9s�E/�׫����?.�x�)Vv�/_AdA��g�@�W=y3��SR��¨��Z3V>˸��]�׆�joY��?e��`��ïx0c���V��}k�^���o��bQ2l���;�{���ʬ=~�y`�Fx�׫���I�i��7q�3X8�Ә��'wLO�z����ydp2�\��_Z� s�4M�eI��ۨ���P�c����E��+�!+��E���� 0G��S�qP�'t���*�s�&t�������LU���n�����
�]��Nm<�����+�yy��YR�q�
�ToΚ�m2(�~��p�b��ͧH"p�3ņ�VOez8r5m�HV#�	��q:��e�:6eE�	f����c�D��ƞ�g��=5\��s\�K�~�ʷ����x��tm��Z=YTx��$]�0?�^�W �"o�Tgi
�}a�x�Q�s��s�ǵC����j����[_����xy�q"rz�7ۍ�[[]L�i=:�4� Хk�{*�I��`e��:�v����f�G��K�����9l��Z~�T��W�O��3!��4�
�N h���C���v���.BkA9�N�>N|0Ք�Kz�>l�C`�n �����Ap�����:��P?�v�*�2�9��~&y�h;VV�s2��N�� V{�d���P���_�%��15�פ�lBƐ�����@|_̌Ss-(��D��<x�ե���C�t�1qfS�;��RcP����7��1�y
npw�K�o���k֔<�Y3���[3�eNq�:d{�G�K*`s�r5�U���^�����{m�`+m���c�5���q����wW��V�)�����1q������q�>�R}�Z\�F��l<u8�Զ �11��v�_���;�oZz���TR�Բ����#�Y��h�V䖙�쪬��8�R��?2��c�D�(�g/�9-@���\㛋��C+2~.���O"�,`9y߭;cC�0I��݆!�1��/�e��8azE��.�D��G�-+�j�ڇi+((��̶ǲ�$������x�k�,Bn�8;�N��Δ|y�z��F�,��AO�u�Y/l�n3�pü�U��q���z��!���;ʡ����Q�u�pd$DA�-�[r�Kݴ|��fg����W/p1�xV<6R(�Z�|�@�om�p� +�N��xG 󏜂��<ž�蛶���~���������� ����d������b���W��q+�+wmaz�K��řcmqF|>���}����&\��������b�~z�1��EO^Xx��)����q�*ڟ�����C�]���[��N�ϟ�d�k?���b�/�u� ������
�R����'�:����q0;��͡�!���li5 �E�EV���=����@���Y��k����7����V��u�� ����J[j�y+B��G�7l[¼oo;�Kʗ���e��*Y}��<�@�@��\�<�������T��C��kh��pgH|������+1{���^:b�����e�ՙ������G?�T��?��G��
K��M����
��xQ�����o�E"k{�?��wp{�.i�?�rw�b�nj���jj~T|]Pp�`^I����Y2���q�'H�������+����i{����O�����[T΢>��������Џm���g{?��ժ>�}��!��ݹ��:�ܛ���`S���D�y��3G�	��'���P�a�O M38�h�l9J;ln�c�ʆ�%�b+��ư��ʤH���-U�[��R-�a��jk�ua5�l�uF�i�Ԝ�`��{05Y]�T�l�)��a@`4�[n9�ΐ���qt�_Ǔe� I �)�������&�{.0��AMʁ�K�r��'q(2+ $�^���.[[[���q"mW/_��	�j�u:�8L*?eY���7>�g����cp��Gi�!�ߕ�?%T�~�N�0���[ =��(��r��V �a���H��Ҥ��re<�:Y	��!����/B�|�[`ܤw���r�ߝ��{�O*;��7V����0�+���_̄k-�0%�[;���R�	,��&�'�uCRF�V���B�o��]�WW��my���m����=�2*���5t��#vo�L���n��?_��ed��f�.D�o�4:}�\�����)�n�w�Ա��^�y�fw�8�_A�)Gϊfnh�G<RUU�kb9���������َx���|8� �BI�?&�E��Ш�����4(l��&�&TWuۥ����`�z��Z�:D���
؍7<9��$����sT
4raa!=�EW�X�������6.��ה�g|�_S=�6��YQ�u���� �y~�V�E[pC��5�^��37�����9<Ţm��*�g�Yc�ƎDEᯮڜF�Y��N��������������Nؗ��9���5������3��V�s9�o�zv���*n�4���@�T%�UI�5�x�C���ʮ��U����on���.�b���]&�	9�B�f�-*˫���0���g���ޛ��MKK(�-p��j����dI`�p�)����\h*\i쳐i�#$��u���Y���e����p�J:�.ב>���
Z�c�eI�)� �I4�a|��nr���%�����JU�dC��Ҷx�������n����qG��[���]B3;��[sG��H�BϊH@�M��R�(��]�a��3�����9Hdߓ�+T�*D���>�Dju)�1o�{�0@,O*�]�u��a����l�:d�U��p�����Mp�����^�՗�N����E��%ЬV���mu?���$Z�X�r5�q�����!Ct�P�`
x�Q���1t�@+6Ю]���#wp���5+b�v���q��}V�G_�^�5]��c�>�20���#�.(>���9�bꊉ�ԩ32�,4W�Ҳ�M�"���l�����Q��;Gkg��RDREu���}SpcM�K�o�¢�h�^��cjj�^�[~(�+t.�S=@���J��.�:|�M����,*�"�Խ���I<-�ע&���qy�E�Z�����t�~{�����%�a0�lܐ��%�F��E闣�����}`q}v��C�:�i,�'��`��Z�{�5h{{h���|H�2(M�/��LnϴŴ�mX�m�j8�"~Q��O����X�������^���\��*�$p�_�x�[��0�Ν|������Syv$wvB��~�`6<B)��8���}6��;̷� V�O�s	���mG|L$��*~[=}�9�T��J_!�ԑ~q,��]�]������CC*�w��n��?�}3�� \rEY����FO���G@#��b�����5�V���w�6d�\�Q�,���A��p�U���'H�/��\�~՗�@¢S��ʏ���W�9�ݲ�ʆ�#���aHՃU���%����]�����&�K��;Q}�-��6 ���H�?8 6 ԭB��������c���UuUU��"���/bf��3_�*��
�8�]�����$M���5���ѳ�|D�^�Μ_x;��3+`�����[��ɏ">wJ�>Rv�-�� B�{�23~{�C(���=��tÌe�<��yg馻����j�Mݴ��i.�(�w-/}�~,.,\�M�P�l��ų��lA_���w���"�x�4���y�>��􀳻���,�h����.J�=G�,n:~;'V<6��̐����Ͽ�-Rns�ɀ(u��p�F�˅g�P��~Yq"�B3�Y�ST��s��� G�A�4d�,����`f�7{wn�ZtS��}k?1^٢�F�?u�D_$�fEyW��V�f�7ql��� �L����� ���D��X/�7S��|e2�G�sq�~��2{�E�a�^��o�h �����?����6���s�WE@�����P�َ�p&c ָ�J�!◴\�R�H�55������e���[��-�5��*r" �%�G���,��蹩V-V����X� ���+�߳)4n0�8�9,(D�P��E5�+��)�^X�4������ �ł ��Yڂܩ�3n��E)�LN&���N���v E�/ӜK� �;�(];S���ڋ��W��CV}�$�}꾍63�����r[hĮ2�0>**��Ҿ/�q/5�rT��\Z�R�D(���f�+g)��&���g��H���'Hi`��%b�2b�@��+F����@g%��&����O�9i)α�}�l��U��ݥ�&<F=�A�\�z��A���T�!;,K���$u���M���?\�o -o���_�r[_7V;�=ƾΧx�4);����������L����*��V^Zڽ�y ������g i�j9ô�����8�A��tէ�1H{��[f,F�-��gn��G��ؐ"ǋ��"��)��nv�Ӣ��3��)����'2�r�a�[���}"\�s�IOOߙ+N��`���$�a� k/τjh�gŘ��]r�.E��wq�ӛ/�#l�k�H��0D��ka�L+w�z.����{�4O]-s�9~��Eg�2!+:�r��?R�L�'F���d��)Y��SF����$ �s��k��M<�3��J���"�	�.r�[1�g�(��>8�L@jxu��~T[2f$K]�zfV�̟:X�q�*��.�>�r��HʿC����jϞb�H/�Pm��	2�೚dʙ��_Ѽ[��/u&����fm/���i����|�r}U�)chϘ�v�D
���w��D�(`ڧb^�꧂�'	�d�V~�gK��h=�=�y�������K�	,.����X�mQ�"J�|Մ�㒖���G盱��\F.O�|j4-��X�e��	�l���h%Ԝ�
H?@��(`s��i��"m�J7"Z(*!�d����a_ɱ�����cq!u�	����8J��79�H�g�Z׀d|�i�8?�;�o%N�~��$�\�X���v�i�y釜����c�'��h%&�I�5E��q�h�bWF��gcc��}���Bc:�-&^M�}����o S{񆓽:�7i��Z�`�;�܌Pv�-����#�i�����<��F�t�ߥ;E��gY4�N��� d�k6��?��xz���;$OU,HfG/4�k��{���0nKz�Kצ��w�3�����m�`vK����cKk���>�����m�ȉ�M�Nf�c6�O��W�Mmoo/��	)�@��	f�-o���u��ϟx{��\��I���x�N~��v?�t��3�	eC����-c/`\��E2��>] Sw �mc^��:�me��piF���ޓ`��?u=����s�VMB�p�=Vڞ�b�bM_3ՎW�O1�K�o���#�v��N�m&�8�	-]���������1_ 4~[X�(���@D�G�/I�o+)��,�Z�V�*)2�d�{�]ׅ-� �XpՊ����r_�l7������K�~�`���O	��'v�YW�+x�,2�'�³�s��3F��m0��.qf�v��E���_��^\9x��͡�bG&��f$ʺ��p��tS��A���X��dd���a�˻�����e���P�� �n�����	�q� ���|�����=��N��vN�Y���� ���s\ �v�7�
��˖�_}�قV|* ���8j�U��|tz$h{I�=k�1�)�?���q��*�*��铼���vVDO��#u�"�L��s��r��7.?Ql�W��*8��ڞVo�U�f{�>����q-]u����%Z�Pd��s������������D߇��]�����E�AN�]�U�O<{�4�UM�����S�9���t��}(�d�	,�+����̫��6�U?�e97"W�<��|usդ،e!�
�q���b�zWB6��k&��y~�RلQU�6����co}�Dt��XO��1����[��pg.���Mz�O�W��Ga��ʉ��W��[��V`��C�biG;����c�i�X���(y;z#d,Uzo��`E_U$WϚ�u+��:��<�y�����ni��a4�q�*��������Ò�f�S��K���Ɉ,E.��6��HI����UT=K_~���#q�ojfb1{�����#d����|�������B{��]E� ��l���ڢJ��:Ķnt��k�}��VcJ��eLW���Qa����Gu����_�csJr��*1Q�E�����(@m���YG��h瀄���¬��==�9��{xl�Z�'K�*9	�X.����"
Mo@��Rn����p/��!9����5:+�0�	��.�Wh9_��4Ԣ��S���J?N련S\���5*mo� 6��z�
$Ƀ+�8D�!X���8:�N.o���x��%�A:�@Ab�j������b�@G�����c�3̈́�٬��һ��<'n������p�2�ZhB��G����3�_^�s�zI���V{����ū���|?�{+�:V�L��ߌ��fK�D4�͑� w
��iنQn��|��pκQa���ٿ�#��i{�~r%����!$M������O��o�R'�����/��`���J={���GZ��/���Oa����
;Z�$�54�����x��Y�E��3D�b;6�K���
�� ��KHC$�[�Ȕޏ��r�k���Mԃ������QAZ]n)~i`6�D�1*=�Lq�(��A����Ӿn�T7�V�tQ��ڽmr��+;*�nw\0�Y��.?�S��y��,ܴ����V��ϻ�̜�L���C�yO���9�sx<g�ؙf���c��h�|�n��Xk�5���(�~
��3����I����{i��{��]<-x���O��ݐ��+Xr�^��z@k�%����d��e�*�n�еC	-Z�q��Z����\l��v����(�)r� k�2�����o2U.�ژ���Q�0|k3�	Qo��p�'�j�om����ϕ�_c���}�;��ݢ8/[�K76\�:�o�\ꊯ�1x=#=�f|��*�v�܊�-�VRJXX���&�w�{D��ApV��+��v�!�Z{ӸG�tb߳�H>����Kaѧ�B�i�Gs_ s��a̅�E��^k���j���*��ݙ�Y3����\���*�7�%�b�3�Ԅ��gPOA����'����L�X%�-�:H�����D5"X4�۳�/��J��w�.T�/hW�q�F�T���+atMӰV)7^�_��G* $#���������{��k�V�P|ޥl:����0UEHC����8zn�/��sj.������2�'e�H�=���6�>.����&�iD���ߖ�f��Q?�J�%lȈi�½������Od�K'E�<:dv-�]��һ�P~b�K����=-M�����E2"0ln�D�{�벒�A�q��K�]���'|27�r�y]��Vd��/ۡ'5�]�����\��IM٧e~׼��v�������y�`A�&��n~�F?���p���x��x�A�j��h�Lɹ��w_��_e�]����v���,����i�N3��w�i�yu|��R�2%�����Cs]��9��נD��XաF��x���,�):C�6?��� Ch��g1	ktB]�����雟A��yE�/�ESI}5�w���� �)gr���ҷ����K��	�ډ�%r\LQŖ:+=��H�JjPɅ�A�Ǿ�@۳��z���u:K�]�q�:`#	ǂ�xf�}K�H<�u��V U��Iْ�e)�ݻV���w؟'&����8�> ��%V^�R8:�>e�l%����"/����#WK�[�Z���O,]���l���23�� ���CA�������|�} ��=�\/�	���1��s������*ZRc(n�"��눝�=5���ѱrqWb�
V��秫�*?��)
�d��O���aI����.�>!,+_gc�a�U�Iz�f�Y�i�z� �5x�7�I��>�>���j�b��+C@\k�?|�ۮ4�[i�*O@zt�0l:~�O��1U��8�/,�/�DEv�!*�g^mw�.M2�mF�h]^�ƗW�T�;�W����
<��cϹ��t��dk�Ir��UR^v';x��h4sH� ����Ut����xU/���3bT�� =R�B�L�������B3�ȝ�(:j�����eѐ"	�ڼ�	{#,��9 �|V!Mo�!�qQ Eo�|�%��^�W��%9<�G>{���HYK����H��x�d�عx��ZR��E`vm"|��L/���a�m���p86�Ƒ2�)s;3�K�I�mV�[\�g%^�Oy ۷��MYih��������%���?	B�����~��V+���68���0�8�8��P,*�����Tٯ�8���P	�'0K���f�y��'�����n ���LN���ɽY����9dD����3��;�{B�R��贃50�F߾�TYW(�34���➟
ӑ+�����;,;�ǭ5�z^a��N=7o�M�p[.=��7ߛ\�|���Z�'T"��F�u�N	��<u}6�QT����?��Ja�7=lFоL��Ʊt��i��[�"�������P��0���N�ZE_��Y'����GR��T�7�n\W���� 6KՀ.8�yă�T�c�ʀr)Rj����~��~�����s��Q~L?���g��b��aKLtw�����1-mn��5�7�Gڞ���}��Qwgv^��No�r��������<�!n:m��]I`ar@v��$m�B�X�,ߚ��� ?����]ב�-K�\�`��^�u��� /���m	X>��m����������������GA� �R)��nP���.i�`(ii�n���b计��3�����u>���;X��p�����u?�sog�`z}�с9x�<�R,�8��ϧ?㟱���tS6����#�W{�W���o:�A;�m�b5(m�e�W�9�M�Q�q3+��YHTS�����VܘnK.�\���WK!����S�����SV��߯:F�fQ���#��C䄇��\��&�AS"Mh������>��t��ts�*�G��-��U� FU1�	7�������>�G!A@���Psl�|��劣�?�e?Қ�y���rg�����������K7w�ɠ�������aH���4��g��a��\&�7-ѴG�qU�Ը[��ݒ�[j�)\*0�5�p|J<������-.�h������^q�����{�tF{'��j�-J�WsM_Xi����N6jl���z&��F��`��?�$��g�o��ϫ����Ղ��$eJ��!��3��C�i�)���ASS��[|�\.p�V!�6����nC�?(�����4�\���N'~룃��h	]�N�g�r�G��\ɍ$nE�Y6����kZ���N���S��>OSb������h��,����pY�,u]��>aI�1�`�f�*�A�����uu�?��������#xLL����8��@�`��^���`�\��9�i>z�ɫ5����,�Nc�A����T��/�����җJkβm*ֹ���q�qҋ ��N�|tf�����X�ʴ�
�g4� _	o�,���o�h_/�l��t����_-v�1���g ��rt,�T)�Lt�؄�|�;�ƌ<�p����������f���A�����/O�^����I;��f�?�����9��Y�a���2��wIR�k��?��!0m�Hd厜�,��g��\*�L3�s �<��&*��o�p�F�g0�p��4S�gFZ;�]���@ȂiWl�C�����ޏ�	 �7U��u]&�>$!�<�w4u�^%aL�o;��py���
�朋	���d�@:���Zc��n�݊L"���oV�v�Afi�|�r��W�����k+6i'4�[�wn7/�à���1�@���#ˊ�`��^�����j𾙿�ĩ}wu&T	bG?�%��Ar�f,��n��D�A^2t�����.����>�����ٲıwcP�l.�(��`��|�V8y�v�*r.q-ȍB¿��=�;�/C\�2X�޽{�S2ϝ���'/)��x��j����y!6!�ѐ�l��a�y�6���[�I�6?�B�q����l�Vx�yx'��ٓ�.��d-�D
z�2���֑�3h����׷>c�/� J�m�07x��o>��+��+X�~����[ڠ��>jG��y�y[��?��D�˷�>���S����M��M����������H���ĠSP|*�}�m�8ԒZ�w1`,�Y�l!��'��4~��T�y洎����;�u�<�� �.�8���i�p��T��ܟ��㡶ϐ�������H	�Y�����ZB ,^��C4�ӟ2ql�z�]-*�j�rSd��HJ{�'�!�r\�v<�ǰ{�Dh~>gE�# ��p�o�A���mI���b#���{Q1�zZ��ΊÑ{�F'�UtJ8]�����ߟ�����N$���/��VUӔ�����9�a���)I\���Ү8V��!EcR�W���b�q*�tw�t�$�$*��V�z�r�N�{ԑ�~l�w�W���b}ܰ"�f���`��_�|*�]h�I:�y��1Sl�Og=�'�M>�=��E}��Si��d~5�.T���?��(.Öv�w��s|�L� <�y�O�+B�@��@���$��~	#�M@�.���z��%���(�9�|�<���R��X�_b�������7�f��aU0@Rk�آ��)�X.�o�0o�>	�|�I���VV�ǚ��Zww��mId�W>A_�2�^��!?ɟ3����U�aģG/��+�ڿe���hn^I\ڣ-,DՇ<�17,}+��Z�1��ʑQ�<�"r�����V�3Y����I�z����Xg-��8�l?`�t�G�U�ɒG���#��b<�
.�NR��JK0�[����S���o��1����f&��BU�6}d�<�Bz�<����j����}�ָ4��x`�\��a�n���?/g߼*W�ǅ���S�92�`�!��Mp�!j�~�$�����F�0���tԣ	���aA@�K�
����%b���@��s˔1&ꟼ�r�/@�:|7��r�~��M����T����YVy�3������/?��C�w�|�g��a���{�xX��GQ��V{l�4/��w�����f1s��g���t��Vs�X�%E|�~t[���1m�k0�>g�3t�h�.6�p�� 9�������� Y qJ�3/���f�1�~b�WW��(>��c�<W ��]dWQ6ջ7�`8}�F�7�Ihd�� ��$�b����]����������jt���g�+�d��}����y��6��Ѿj�g�c�B�jP�S�U�Gud. �"d�}!̳$
 ��eSZ[l[�Ԑ�I���D��-�,�O@�"�D�\`�\��������ޙrh�膼#^\R�Y<V9Zٟ�ݻi�'�ŗ��7���K�`�?����v�ȉr8�S���R
0��Y�U�M��rB�%n��N��/�2�w�o�0�s���� J����m�{��w�,�v^�ir�O>6,���b����µU����A�E��"�Ky�9A�^�nvvۨ�	���^��4Nd23����ג���/U`��'�t��b<���{S<kS�R@�	�tu�}�8�8F�������Ǳ�6��TC��D6�M����Ӻy���h�����{*������ϴ]���#[_u�8�r|]������~�mc�͋�<���{��^'��p�.B ���WXLtX���dg6 �H�����q�C.{���˿��>?J��x�!%�6~�?�w��|����M%�,m���2��y�V4��rlU/j�� �����z3˫Xm�?NFl�\�������j��*7.��$�+w���;����aJ�[�k/=�fn������0���b��pV_�Y]nߘ �q1���0�X	fDZhQ��n���:�T&�i_�Ӡ/��h=X�vÐ���K,�]�Iʁ:�/��P����˷���ru��t��S)��g���o���20q_
䘹8�����y�z����Du�Ju�a2Ӛ-�G���u�§�.�q'�%�>	٥��K�3E��&���ݷcG�!���J�"����I��;���fX��;¹����gp�������D��nӾ�E�h�@�z�����HX&�̄��% z�� ���xpgz-�3���YW�(Z}_�%v�엗>��]sJ��w���m�q��U���.F��\�\�δo	��<�����?��ڽ�X�6_�ծ��ɷ�s���>����U�}%vDAC!~D�՟�b����
yE t�P��vO��������.U��S�lU?�+SA�`�F�\=2�,+<XBN��C�쪡����ϲ�,��δ�,�w�)�5x�3h�w9v�7�	ַ�Ɇ��D�#K�h#sX��t;�fO�F��M�Wf�te��+S�L�F���n��М�ԾMx> K�/��i��u�������w����3�W����//���1���B�5��:��^Oz�\���%����h�D7vzy���>�88p��A^��g�Xu�TJ �؄���#ݠ\�#:|�z�Y�PI��.�q5��nY�bǟ}mϔ8��tOprL����U�;1�����w*:�{��*�,�7�K���qZ2��	���:�p><V�s�R�O�Ж�ղ�l� �?�b<CO�l~�z6=~)������S�G��3��J�W��8{>SN6+\y*�p�@n��-SV���)�F��.��"��Z~����-������k�0�MX(΄��ne����iL̐����m��Y���\���#&+= /Gk�ȫ��u�PD�3�s��g�_v���/9KKҰ�K�g�ś��N]��r��<�Amgx�:o�S\-�����&����;�hE@�U;�G#X�6O��`���Dz�K*R�픭�������++,`��9�oq�Nv>[�(5��A����Q�����D��?y���yQ�5�,�o��i�J�������N?�}���"arw��T��є�`�q�Fo)U�hd�o�eǠ��{��Wr�����?r<�.Hcb}���*��I�%cg�(Eg�:8&B<y����ݛ�9�Շ�z��	<�[*M�za��Uz-����/��<��?��)\�.HB�I�nX/D����3.�jOt�B����M/�ԗ@�5���8���k�w<[�+���o���r���s���@�'���+����:�~aF���D��NE󺈙d�N:.)��pI�jl��H���(�ٍO[����l+J���sY�d�����.���eU�g�/ֹ}������Ger��T�����3��`#H������A�g�>%�s��͓)waXD;_��,I+n8�����D*��PY�1�c���;I"��4�򳻟,������3������Nl;��@_��I��+����Y�3�f�8��O���f�6�g_�+{zH��l����܅�����a5#Uğ�诐�qO�)�V甕�;Mşʩ��x�v|󊫢��#&D7�ԩq�nGt�pS���%��wz�a�Pj	���~�?���R$�L�������q�m�D�A�R���R��E�ugot���[ɋ�+ؘ��DF]���K������n]��ܛ")#�����I�
zR�wW�%��/ֽ}�Dl���V���U
"Ɏ�H>KC�G�v�8	�I�_�ӿpS����>�]P� �i��gM/.�������(~aJĽR[�_t9�������&j����?rl�}D��&��Q�z�����Ż�m?Y����/�Xm?��E6�]�[�W�	�K(��}�����{�tt��a&!�cs����2��P��QO}'��m�XK@t�]�T�����O�D�R~�h	��r�{e�d�Ս_��P�^P ��>�D�o#�O:�h��"�
�
�DA�닀�a)0[{4����t��R&g�8�l�k��1�!b�j�&�� n����	&��DQ!�db�O_�B�?��g��~h�|���ռ�9x��Ӵ�	�x{!�Y�%�ݬV�%�i�kh_#�+ԝF��U ,���&=��4��=�׸�U����s��?���u�ꎙj[b�(a�˯ѱ4 �"��R��Q���V:��/%�5��B��6���R(�����j�u������{0���-�����j���'� �ۦ/��S��ؚ���&Qz�Dur�EG=[��\vJ8?�Y�jD��~�w�u}��G���qJ��� ջ�E2~#}��gM��.���E\�����ֈ���'*���\�\�x.NR�v?��ܩ���.^ ̯}�^H�A^��N�O3����IX-���M�f�X���~�^)ic�H�5������ꅑ|�KO�[.�(/�I�H�8l�s����k:�D��ӡTD�⹣,]��Ey�AP�A�W��I���?3�:�3��U��y��p���L/Duه��K[96�1oŇ�9V��(��|�fa0LN�t"���v�ua��BV�#�IgjbDH�!!ci�b�Ȉ�FJ�<!�7��.���@�5}8D�R��`"�p��GL�5@�ɑ7k���KaZ�q�,��Tn��P(5��l����)sC���Tc��=<[_�3�$�Q��$z���c��q�S��Ð�w��͏!�I������%TU]��-�}�]CAy�j�;?H�6Z}�Z=N������zP{���OD|X���r����1[�[����ؼ�x<.�~�Z����s�*	�=D%b&?*a��~���q5ޑ,R	1�x��F[P���vE	=�0���Ȓ���Г�?��-�[��.��+$�z���_�����
��N�\
��O.-24<J|�J�|��|�H���܄�8v��Äf��+�y����B��6V���pO�*��i%��)¼�th�1~5��~#���z��ms� �5�atO��^�����K�����|[��C�h�:/��f�:���TZ�r\���V���ӎWH�hk�>Z�࿭��}<�ڭ���Ye���2O�>!�wQ�i�i_�)U�B?檨(�O���tߧ�4T��E�Z�HjN�%C�ݒ�f5����6q6wi�E�O�d�Q�[��#�,,V�D��=�u3�WCJџy6�Gm��53V��<�2�y%�sH&�{������{��l�;���3�GYn��H���'��y:6�,!�z�{5�|���s;3L���OF��J�o&c��~٣.d�+���Gµ�I�@��/k�x_�Oq���;����ℼ�����Y���|��W,�x"�\J!`:�X埍7Ӽ!QX��HU���wةČ�e�CJ\�	��;�ϑD���&(���'iH _��&9�h�i�{�\Ba�ɥQ?����ʰ�6��qu_�'lLV��%BQ#5I�$^:I�%��b���W���x"wq�[�om���K�5�_\s�p�';^�|4/����Q
d��s7��@���3���������K�B��`;v�VG�#��Q�W��K I8Yn�#XPɬ_��N� �[�eΦ�,~���|+�YG�F> �r�c��
Y�`�J��"l,_��(9F��ee+K�իc��q�;�����}5�����|��r�5}Yk�-�R�o�]q��,&V?�*k]����� �^�G��(�d���a�Vrڝ��#,Ϧ*XUB�2���������W�g�K�u��~C�\�
if
�Kj�~F����Z��>�s�}�|��.3�@��|)L��$u��W[B�k�ŗ�M�՚��'��X�L"�N�x+',%5�a�*D��t�y���,TR�ʟ7G�i���S;��Pqp�F��p���5|����4�����]�Z��{�k�'��Ԇ>�}�s/��y�
).ׅ��p�c������:�y4y1�X�_ǌ�i���>+)�"@Xs�Ty��͟��R�ECn�Biǒ !^�kq�ѥ���J"���:�#�)[&g4������ �Vo<��|��rvm��s���f�����:0_F�ť����j�V��0z8!�l�yP��0B��y��
j��R ����q£o��"͜����Ř�D!+sX~j�q���kt��a)%���D�⮫�P����b	�q@�!�kB�5�"ʼ��P�rr�lqB7���<v��>���,2�œ�/}ᢛ�=�|�G9���Kv��q�E8A�%�I�4���V�!fS�2�^�=$��c��#<�8������lW�lY���_xL�Q��rs����a�<c��ԟp&Q��Sz���t�ۭK�yG^rz-��U_����-4k
"~'�T5��+Ǧ��I	%xu���=�j����VpKo�p]����}�����B���0�����T�����BX�XR~1�cF�K����G��A{�d*?�c��>�Uv'5�����Ӓ�k��.q˳���.���G.!�UN�k$����JA8zRg�|�l�B�*�v�cLh+1�����%�o¾�H��5+��2x�̭"|
#Q�������>��j����f*a#S�r(�&�1�nw%t{`�ʗKj�� �v9���K��Ce�&���3?�-?��:��+��� :[a�܊}hJ|��
W����{��R�����NB_��!�e��D���}�f2����8Շ�VZ�V�+�z,�A�R�n�"�TB�Dw��������e t��;�Մ�����(����<�
�R�|�����G�bS< ��Ƥ�t��\����up��T���x�v���ܢmB%�@yݒ���oxN"9g�̺�Vc-�نʢ�{!^L�ۃ@S5}i�i�ߴ]�M$!H��#��_U׬�\��(���z�/��ï�X�D�Z p%��F!;c\[Ŗp	�H�ȭE��QJ��A~���p�灬ڼ��+��Ip�[� (�M�����@gx�1�{�&�濧�M-��w���:�V��$��s0�6�{��S���0.����7?��y~8��1.�  �&ݏ�����7eb�X
P��n}��~�jb��`���퓞�ƫRB�·<�(��;�@�����T���;���V���4��O�f�nX�W��~�!��Vytx���8�#x�� ��(g��.S\��{L�}���M��:��~����d+�NK�0�
B%������U�ч�l����5�Ϳ�0�z]l�,��h��Te5���]]�E|!	ց��X��Z��k]��XNN-ry�ż3S�������QY1�6�raα=�%�ki~W�v�X��X�ծ䋹(���E��������sn%IY�"SY�q�jP<�|z�h�0���ӑ�)HiN�m���LKR���R����՞���=� �V΋n=6�mmw8��Qۣ޽S�ɝ Ą
�������0��x	5������|Xk��zP������ir�jS��r���=�-�����&�It�@�����b�5M�I궖�������?b�Y��c!-�����#���e�u��]dNc��\$�v�y�]ȥ_j����Jn��J�/��o<e�<��&�9��F���n)aR*���a[�G�Ѭd��b��ǢL�	"<:�!�{���ے���:���9��������Y�J6���<B\��[I�O��G�0���o8o4Xm��uk��z�m��T>;��X�u����z��Z-Z��I�{����&U��߭�R⏽��٬�P�~���~��פYr˶f��`T�TF�&���=$t��xҏ�,�I��s#�
i.k����@�Oo�����w��d���Jh;A'}޽iU�"�N�����?ۉʋ4Jca���܎X���7o^湍*[�����!�f�.ٔr��iw��	Tu����NTr���T�}�q�3S�:��a�>z�v�0sh�i�AC�R��:�/޻�kw�IxqW�}1�)�T��#��xՍ��I+��x���8.��h�-�`�D_2ʉPJ�B@o��Q�j��B�J�����Wy��ȼI*�b�v^=<���+\���̜΄g���놿3�@.ҏ|�j
S�JE[w~����*m�-�=�m�U/<X�8	��0����Fo���)��a� 7lf��2�j�/%��7t�z�#m�n�.;JF5�a�Ys��B��]FJ�ΧS\l<�j�Cd�.�kj�)�R)xi�bκP9h�|H{x���J������{�(�'&r^��(����6�6��[�!@=Kh��]N_�����#��ٷ/gM�'�q�E1'����]"%�������|&�.���;��<D����V�|b� m�k�eKѦ�C�}���p��xu�1���*iQ�/n��Hg��[_�,.��r_g/|��	�]W�xz΀����{d �n>��1��\�1 `�� ���Ui��@����|3����W;�}��v���D�1k//Q���Q/���o1�6GNr�ȴ]��b"�$u7ϣ�F�M�e���AFғ=�zz5�����!�	"o�ٜi&�G����z�1T��H�X���ao�ڗ�]���ҶqD���N6���G0����&*�	��j��㾺{����T=�o��[H����8���cá�ԙt���ՖK�`�o'��WO���//�ը�]�T���������l�!N�[F}*�<lĴ�c�.'>A'�B1�ѷJ�k���g�[��]es��tp�:4��X �B~a E��m�b+��ϥ�.yI	�F^���F�lLT
G� ����<�υ��#�ccl:�C����z�Aߋs!گ�Oϲ�m�q���"i������	 �|
m��X�!��і���U���6�	Vs���-!�/���>��/=-��lNj������XQ	.�C�,���Y��ND�-N��x�l��Ɉ g���+��-�?�/s$�l�]�U���m=zi��7��5��xw��4��YC�P���Y��T���%`�=�G�ˇ��=��_���>��28�O#l�� :�׬Zt�H��B��Z:����dip�"�Ash8�&E��5�L�R��\pq3�����C f~�4�qJ )�m_Px���H���,��ǞL�q�-Kw)�ץc�r'g�M����6�¬3bpJL��u��� qNe.�A�ao^1}5���ҁ���}�1��e�/���TZ�����-��>u����k���-�x�1�XK��߼e����S�ٛ7o΄J�������0|m惲^�N.�_�=����8���:�	XIK�Ҳ�7E�����/�b�[�Z���O6���m�r]T�y�~����\T^M4��U̖�9��o��8�_��:������v�jBg{Xb=F��?�nb#H 0�Y����4����:�_����������E>�~Ja�༹�,�ո�����@��;"g���t��R�d���VU��X�]���N*����]�Yj��-���׏1�pF��Gqs�1L����7v�v]Ce��j|=='�00�����|D�=��66�ߓ����`�V__��;m��͛o�`p̢pB7��ﱕ�ʥ��6��G���У_�������S�[�hiy*�~HIisshp�#�����?)i�+28�_n@sb���U���ӕR;�Ð���cu�k�x�x>x�`!�޳j�:x�l`�a>V��cz���vN?؊M�
�5���	F?ea�.L�ѱ赸x��3W�bn�àkU���Y���Ϲ��Ud��p;X����d�_�"�J�6'�g15��e��,����Tw8�5ٜɳ*Y��I����424�agW042�ea�T�,�� �:���<SQS3SUR
���N��y��_���I	�/�Ɯ�(�t}ww�J���&gn;Tݧ��>�=���Q`�5n	y���l2غ����ij��Q5�6��כ/��ӿ��j:<ż֏��tX1�dj�'CK�CG�.�j*3�z�]8!jGɵ��؍�u������X-EI*嚅���\ď��ɾ�Kd���T��x@-�37���64'�t`������+U�����g���7�'�U����Ldff��4G_a 0==o����Xjhh��(�!�n�dc���F��z��pڇ*:����?�mlf&-%�{e�Bp�=�7���h��V��@�*`g�~�E�����
�5p���FM[�����e��S��R,����uM4p����	);Dh�s*]�ls�������b��Kl�pv#6FL��� ���899w���/����<��vڣ��+�ܥ���+��C

樨(�t�u\�W="n����{
C�X�*���8��?ߐV��x�C��yO���Wy����d ])9=]J.�� be[�
�~��i�:�`Ķ��K���9g�����
,��1�9�����ʬWNj|"��:�6�Zl���{J��3
+ڎӿ��b� 6 1000��7h�F�X�6J'�=28h������C/Z��fc}�*���5�B1�
Y̔��g$솟59P(���@V|<%�M|�{��/ׇR<�|�x2�����N:סd�`�]E�iz�z��I{G'�x�����t���0;�ѻ�v��
xo�-��}�U�i��#)((X�Ї��n_k�V�S6, �.~�����ͭ<��Z$���FMF�a-��o����vkw7OCOk�s�D�������Ӷ�����PK�����Q� ��߿�8�}��C\���Xg���F+���]z$��Er�h��/�JJJ�:�, ��q����>i�q�e�kmxer��79�z�Lb�;�˽YX`X�Qs4�H�����3��;@ӏppp^����q?�ZX0u�>�����r�?���v��N �V\�����ipPg�Ty"8�$��`��I HBB�5U�������RJK�/~'�.� ��Bw=K��46�&r+����kHU���$����_�...�p��D�n����[?�����U�ȬX��͡�:�������
W'\�p;]��D�F)��P���e:$�U:��� ��l��n<��Z�����Vknu�D�).�p�ܭk&�Y����cF���:�p�W_!�QsQM.�� @4�O�Ǳc�����Sw�{�_M�}�&D��4j,zm�B���uŵ��B-3�ř�����?G�;eDя�xՐ��y��"^6�%�$�z 1�s��
���0�;�8ٗ�� ����g5kU��U^i�I��j�����:���d�c��x-EB���`r>EX0�|���)�	69O���X�w���5�v�4���t2?EQ_Ԧ����V�<�O�}��J�.��MW�^KR}����'��L��4r� �-�I�8����VU���% ���SLb��X`H8$���&&&�g�x@�Y�Ѧ΀�ʴY"�>а�ȡjZ)`Ff�FV6����)hԠ�H�0)1��ǎ����l[�x�\V����kP����U�������AT"67�az=�>��|�Qۮ+46�I��?������Ƌ]q}==������ТxA�@v��O�vhD���8)0��Z����,�H ��[��U�bQ���o�N-	`���T9��D�`w��~s�6/�j��3s��q]���ʒq�!��r�� `T���Ond�an#v/v���(���:9�8�
��!eb��V�a�xS���D	{@]�kΏW��X�5�o�pW�iE�7(����N3nW�l��UTh�Y0[x������ܠhΜ�-�ˏW2��&#u*���.$�k��)�8�C��_�	������0"�{* F����{<����D�U�%�>���z�)�~��D�y-H�W�"j���Z
�bF�؞�W�l��;���t�St����Dڏ� ������v�JRvû��D�	����<��=�8D__��\���T���3��&@���A#ʦp�o8Q隵�o�{7�H���1�I��������U[�lNa~l�%��e����k�����?�n��}��F��1�� ��"��a9�D�m��0A��]+R����5,���D>ODَo��Y��ݱ1��HH`UJ�y���\4������P� Q�O���G��<.4�6m���,��D"�C��iQ�D�\i�?����_�<EkԞc<�c���1�RQ��]v�Iq��u1@��?	xׄ��Q���n�d�UQ	�6�Z�������Tiu�������M���V�!s->xܷ�{��j�#������; �k�s('�tW:���ޠ�;��T�: �����-|n��{����+*��=0�Zz~�B�oƾ�V^1�att���ȟ���ε�v��բ� %�%%�xs$~����Ѩ��&�P���©�S� ��V���&@�o�ݢ��_w� ;����@e�N>��8�ޔ��1w��7t{�t�e1�,tt,Շ����h�ȑ��R�$'�Z�V�			a\k��	 �(�c
���H� tea���I%�;"<��F)�c9ڱ��\P���|�^DD��J����||,��/���e��}2���<Vb����J�s���
N�\�0�K����G�h���}�O�T���o߰/g	,����'�-��:,t|��uD���¶��بfD�_\��\kΎ��˗ƣE桑��h��P8*#!l�Z��v/�c
����555և��i��M��C�p��=`��[���5^�iX�2sS@o�y?��@B⍓�ܾu��U}h�Et]�	���␉���t�UXX���)4n=dHΓ��`�w�=��y�fvG���};̗7��ù��T�]�#sKK|Ln`��m*I8L2ʲ�)�U%%%�X9��  ��V��������)8��_�~M�>�]Rn�	^q�C�FDHa���!@ȅ1�ng�8�H�	kl<<��h�QQ���<�+g�Q*��T6�����YB���꼷ͣ��7��a�IAK��l1�O�|dD䩡�&"Ȍ/�� J�hbR�襝������+c�ܫ�T`�%�x#�h��4�>�ՃT�3)���M��" BE��ӵ������}������ER�y�D��ʨED�"�y%㙪ي�5��9��v����0bd�
c��K���h�>�ou�ILJ����yA_F/���kN&AX��8r?IN�b��#�e<�!BNF���5��pL�Н���5,uUɵjb�F�n�f��L#r��'�c�@
��ng�VS���냯�d� M*� ���46@�_ii�U���	����tFo��Z+X�1��2#p���{�Af�ܢ���|AꎎE�=�I�rm��H��k�x���,��$#�Y#[89���|��Sc^Y
����s��m7>����NΫ#�W}�s(�7�д] �g�N`�m�ֶ��l�Ґ�� -z-!ц�0lALs۲c����G�a�5���P�(��AR��C����9>?��*s�Eu�}ݹ�<(y�0X�͛oJx��1���ܪ�����R�z�PYX	Z�
�K����n[�������J���G�2��pZ�ޮ ����%p&��/6��ms���	ևO�X�_��Fj?��c�� "9??���������f@��9��H>��ʫA�����;V�64��TPP� ��������<���S��Y���N="$�C]9����.���蔪_������cU��=_�����g'���g�[�߈�7����Z������<�b����*G���A+*�>| ����6
?~l�0�j<
=K��B��K�ѻm�ғ-��z��I������;( �w{|���ZE��������Y�*^�v,Cu��G��`i�wn�^�J@��@��J]=�o�L�����y���bF�a�;��i���g�Y3*��7ؕ���;�;��}��ri9\YY�/.*����\��I�'����|����@�p�c�,��l�ϟ?-WA�^r������w�FF�+�5f::X��􅟼��$��W�Ug� �[3M��B��#Y�_|UTA������l�E�Woq�J(yEz}_L�ҍ����@������1�R�������-;׬��I��S1=L�G�-����S`0ع� joA���M+E��������W�%�Z $�
�Y��~(#+q&�etlt�|iϭh�5�6�lU)#��[�ŋ�~�V��װcg{�'0�D�ԓ)t���O!�=^ �^'��իlK�g�A�+�^:��8T%{�8"���"+�ϟ?�7�`P�Qk��-��k{m�U��&G�2�=��ތP���jϭj���Yew�B��^�}�|�2 :@x��7�A�䌔���'o�w;��F
���_(HJ�䖔8�988Lﭖ޹�i,�jzWO��g�e�X���	i����Ы�0���L����cqr�STi?6Uu�T��ĜXXX�<��x�l�z��������?���ܳ�s��ʃ��}��"h@Jg�N�9�d�D[zf&d���%�cn��&g�{��Ip]�����0AF&DY�Qwt�p��uʋ�[���O��M��U�yII	=���!��:$㰍����ޝ��A
���ϙ�d:c轎��dd�e�Î����$�
de�҄���?P��;%�0T�"���Z9��/��:�·�BCCm����	݋���a�|���w��F����E�d=�����z����J]�
�,,�f�HA�ּ����z�/gS����?�lv �����T'0xupp$YBk@w��ګfkZ�gB�`�VF�����Z=Oo��~1t5��4�����,�E�8��t�O��������VG��^��Z���������W�J�}-���A�V��4ڦ]�$����,��ŧ�777��@"Ck8ϠA�H2,8�qK��7�zt� X+�^p��h�^_REE�9 ��,}��$�7]�1�ԡ��Q�PM]L��#X*d�^���鎢V���}`UBP;�Y����Ij������2͘%E�Y�Y�Ho�8��L?��@H0���6b�h� ����I1a���E�]�y���Y�d핑����+޽{�}N���=�ˎ�=%�պ=5�`��UZc�>r#&Ȭxl�-y�G_����{V�.X�_��K��6ZZZ�---�/��V9��󘭩���v` ʥ
��� ��a�/0i"k� ��1pK7���}ӐA�	A�����%10+q``��x�k�h�q��,ݪ�_��ek�"Ka�cd�� 7��0��g8/�pX��W�E��,���`3Y���Y$�32�U����
!�n�w�gzڊ�����NŘQ��v;|�HG��n�B?���^)|hh�ĩ�B�jh ��]�&�LLL��LMY�+�Ŝ��hud��D^'�ĸ�*O��;�,ﻵoL�;.��a��X�%�0��%|��,���-ϔC����������#�e�uf(0 $��N�3T�0N)r�<_�j��sǉ��JM�z~�|\��z�6��a�M���iwm�v�A������J�x>�ǅG;�'���������iiiXМ�w�EO�(�ts���������E��3[�������@[�k [���`��Ij�>���nki������?t5dO�Q3�5z��Ђ�@�<|��V��s�?R`�~3���"r��5�����|�VN'��X_K�>{�<~�?p(Ü	lB ����S����3�'�ں��I}S� V���O�n�������������sʚv�|(������{f��M1! UN0����v��.�$	����Y:���yU��'���+f3����q7�C-���c���J4E��O�jNrqkk�����<I[�i
�j�wj��� ��|�C�z�<\"��z����}ɹ�ۑ5�= j�2=��o\���n<t5?�]����	�hFfFF��XZ��xT���"��Ë_���'�����[� ��w�hw��S���bސ�?O\=����tß����D-G��V�d�(o<w�v�����u�����?}FW�b1����*�����V���������D�#^�|�B��xW�����_^&��-$4�i9��w�ܡ�%�L��њ��L)��/��;�����LB����#{]����*YI%#���ޣ̒��l
2.��<{�^�O����'��s��<���~���ݼ�a��{M��+C�i������x�s�`����oj�ꎨ?x��
Ҡ;ao��R���<���1�G�5�*�����^e�4�a��##F�h��r��&r66y?DuW�.[e�*�?��=,4o�{�W�js�0L����������u?x��3l V�}��"��<p���_��G�����YKDŅ|��m��5�t	��DqC�O�c�"z`�CWM��r`�NeE������k����U�C��vf1�j���:}c���h�#�4���ni��Hele\�f�� �^0::Z���^��.����2� bۮ���՛��Jmo�؁��cu�G��(A�9c,�������"��>��w���{]pn�zE�*��e��ȵ�J��8_�/�T��G��E��7���)z�۳��l5N���I@������O�����Zv�oH�V#�P�Y�z���>}D�����FA��Ŧ�(�XmB	lbbX�����/c����ϟ�����6�߁���p�w�5R�!�tMQI��]�r��V��G��j�������]fNNN�\6����t�Fm|4giiɞӸ������j����+i��7r����|��������`�`~�d�Q�-�A+�Գ2��Nu�EVm&�l�Ӌ�,}�ߣ�� �d4 ����1I$�aM����yX�r���ߚ�US^TT��-�x�]m�
����Mƴ�-�i��`��==�����ĳ|��%�>; ���m�Dz�{g�/�uA8?b�<_ϖ���,7E�$���j�Ye�ĳLT�c��Z�Yi�}i�8E���o�%鵦�#�9�:�w
��۞ԌȤ�C�H��]�L������n>n��삂����#�(����#S>*�kWlF�����o�n���A{ͧ�{�[$�[
6K���K>߇�nrp O�ΐ|Z��O�U�D����E�p��[���g�t�cb���~}u����v�b�	�ӑ�/��eff�G���]�y�@�%���	~�뗀Q���]s*0,1W�(�G��G�T�..6<���4�懖����E�j7F�2+��!��)uuG����8@B��{o�O�X^Y��t]`�EĢ�����Ҟ,V�pֈ+� 
>rQ��s�h8�p8Vv'��a�l�yYӕM %Qp�zk{@M�ݽ���:##������K��}��xR�4y�Y@���6��mD�ܹ�C����D���C�s�m������ѣY&�Ѧ��-���|��fFO>H�\1�PM`�=�[ �c>�������s�]����xE��#���w-KKK�:ٔ+��H�I5)�}y�����'k��Z�7Ř����쨁��Gy�9�\�����o��'g�WQ��1kFd9x={�����t*�{���-F�wvu���C�<Ěb*�R���;��[�����ֶ���cXƓF��ֳ0[ (ob��!%Yc:-^)�ǻ��ۯ�,�F�ؘ|}�&���id�{��n�hՁ�{B7��`��CD@@o��z�Z��tA����~��~O�>�������WJ�;yƃ6�"y}�D8��d����ѭ0S罍Y%A��K��- �T9<B��������Y���[lo.�w^L�w�#����4���nz$rF�/�=��W\58�uU��3�ǲq�ʏȣ����n����kk��4��X����p�~�U_jw]]�i�t��|'�FX����;�2����{|q��v�l,qZ��̷�4�-{Q7O9�O��h��	%���?8z�����zO�Y7<���F{��N���0b`�rL]E~�U�jSPe�G�����Wj�͎�^N�N5x遼��<�g��c�%hz�e�/��g|߰�%r =a�
tMC�\�q�ݤ�׵�m>3�2���Lb+/�����^�� 1�nU��X�+k�E�'qn�nR����-@��z=p�����o��ѿ;}9e��%&#'���Jq��}.�QI���\]�I�G!����jo/g&Q6Nsc7	o��Z �V��!fO i>x������4�ɸfۓ*�ؕ9cm�t���`��ZV.m�����ՖV2;-(�t�C��Xl=��_9�륥�ڭ��unn�Y�Xb�C���í/-���Ή� 3����W4M�èt��6O_{-��e[ػ�t2�3��P�C}j�@0G�lo/)R�������F3IO�Z�D"����X��9YYo���c7+������"��U��7���6�PRVQц;P�#4Aԋ�¾wuE��w��!{��?_�,�v�mZ�������`���w��Y<��,���v�W��3t�/,�~�l����_I�E���g�q6>��I��8����Y��W�["	OmyWŃ���"��a��mm<�����A��E'm�$�a�**��i��n�X`[�n3iW��$:�	w��e
�ɇ��Bu*l,,�￡�u�Y�1�k:�p�*��+b:6 �ߙ"Ĝ�!!3x)��C�vߢ]hx�E�0"��a�տc�?AVN�s�/�u�W[Oo��u#{S�c���̯=��/2"""7bI$�䬝fkv��6222�ː�-�f��4ӱ�N�H�J�JGu�\85�z�a� �ҩ�z��;g�Ϸƭ���i6�ߤ�Qүa��p��f��^������Ӯ�� ��puu5�_�3���k��/�����A��g�!�th�N]��7�_ A��^�w�&j�����0���h��[P���N�蟅F��SF��_�_^�Koh0~ůwF>�e,�pzpI�Q��Z+�x��-NN�Tٜ��ʖ�[6 ��Z���&�q''8�TFv`ųO�Xbj�qI��ڛ��U`�O�#�l�ܣP@^-�M�]�a^�:&׮K	ș�
h�<W��d7�}J�����z��Ɖ��lm�-�"B�
"L�O|��+t �������ʙZ�$����{N���DA��v?�,W��0��8�-/����g_�6��{!�xK�y9�$�:���#$"$��X���g��j�(��W��+�����be���캎�8	{xd� -9���[7ξ�y\;��/�1UC[[���������67��V���q�C��o�Xx�i�¯���! ogW ��q��'7!;�+B�G{Z8�� M1S������Y��,�����?:5�W���Xi>��s}h;��7��1=�B��ԙ��<9�@�[m)܆cQ���2�ETUR�ư�&�:��ָ�[�x�gJ-aa}^^ޅ�r�Ĩ74Zl������Q�:؁?5_-��%���Q�!�d�$�z�� N3M8,��w�D]XX����9���?e�ζL�{��QPV.C~�j=n&��<��{��N���K}��5�ll�w���@��6+�j�� ��ݡ��CV�5v7�B�ϟ?�Cg�K�`�o�L�SR>�>'gj�j���w�����'�]B�מ>}Z�]�Y9�c('��2�!G�^��B�;�|��y���]w�ND+/��t�!p���p_����Suf�_I@�����|��X�w�:Ԥ|��)?�I�vĳ~J�D
��<8�CA���5r�<k���ݕn_�9qgQ�3�F���z[0؀]��Lu x���eaSF�=E��?��a�0W�l��.Mu�"]�aD{�sk(�d��$;�S�Yq��#M���ʹz�01I�e �h��D}hx��\L�����K;��?e ����{}��r��ݻ_z����f ���ݸR#��a�#�����:\BP�4s³Be_�^��$..Ώza�G!8�2���i&�TJP1٭�ش��A�}��tO��ڞ_��W\qng����R�S^	/��s	�G��	�eМo��Z��O��q���s*�t�Σ��r��X"JCS������tVe`�*�D�h=bdg�Q��:>00p�Çb&�\D�KJxw�IEA�p^������W�3�{-y�-26��s���R������xb1ܨ�<�q�h�������� ��l{��'����gm�>_E�I5sQ��"���/C8�ee.�J�o+c�)��{��*���.=�{�؈#�}��ʣ~��:��"�aaTW1KJ��P�����uV(EE���m+3�h�<HC��##~@�1�r���8%9� ,?`�37�A޾��txTVVvB��7Ӵ^�G[?}�Z�\bƮ�Nw��V��=����+�9���;���� D��m5V�[��w嬈%��!<�y�zÁ2n��bSR����$O�{Lu�280����Ʌi_|���D��Y-ٵ&x�����~����c
����^����seWUP �����R�Ӗx�ik(���}�~vO�����:(hk��/q�o>'�x��Q�ռ�w���N R��L�kq|A�"�1�k�eebW((�;��Z���}��+�B��]��YX�4�k _��[�k{u��x���\|�����,�T��H��JS��c�F�>��|�ҝfm�库��=i*f�b�\d���'k�ڴ�n���4�,GzE��8��+������A7����?��c�I�o<�h��K��J)�h��7K�2�(g�j�҇ŰV��3h�QD:@�����BE��t�q�e	����l�>��,8�!�w�_2J8(���ښd��r:�:Ý��__�y�_� ����G�^k��^<�a� !�d "�gz���:""��H�����#a�Upv[PB���Ug4�(đ��e�PA�[�����ϙ�J������$��6!���Bᢂ�?�6�R�K��pjV�� �]ؘmƚ���`�mSRR0D������C
��<~�Ⱥ:1���E�$|��������t)������+`.h�x'P\f���ê�g}n�ݓ�ffe��XH]�+5����4t���		��ʛN��q-K�P�Eh���������ϟ�&A��LSxk�����+���&��:��)3nQ�!����C6���J$��ߞa�GJJ
���G0P՞��PA� a��ZR���8�?'���������Ϥ�Z�u��'�d�[�L��̔�}TX��A9����x�{-ؿ6���EQK�^��Tb\�g-T��b���)�u?��(�����e9R������'�F��_��b���k��@.������;�~'[I���~��d3�<�d�8p� �π_cye ����>>�<��m�IW�4��"�����F^��S�&��ooCC	�_$V�~SU���J�)��F5TT�� �Ղ��z�t�yJ�Ǩ���8&���{�� >��&C�J�w�ޙ��YX�_�a ���y0ikk;͛��J�`��w¾1_'�X�wH���R\�X@yhA���554~��o�8|������M\\���.�C��P������i2�bqǳ֮~gxz��ϓZ���%+8��Ԉ`e����O�XtL��$)����1ɞ���|���yG_��Cgr>w��l�u��^]<����󳳣:j�>1:����g��u�\�c�y��h\���4p_��6y B�3v ���Y��ӋDzG@E� [�A7����W��t��h� a���[�cf^^@'[]�^����T��O�r^�,@��K�	�,������+�=�OJ��ںF�Ν-�����͌\\��iX�r��E��Oݺ�ѭ��<5���+'�c{
��ޑ5ݻw��o��L������n�6����o�A:�����~�*/	��]�߳��g��v<�@_��w'u��6�
P�
�L3v� S�hh�
23����������A��GB�'���I�Ƹ�J���JI�{���x�����	�]T������:.��֦�r*�KZ�44�k��uC�N��S�+� X�wAm�|�;_��e�_�Z�eJJ�^���qP3�1����˖�Vi�z8�tt��K�������U�akY]�8 ��6]zGx��i%�S1䄞�w<��BKFA1���M�o�9�444n���}�7���������2�r^��'ɸ��1�-mm'�^zbb�
@o��m7r6]��=�K�55��e�nnYٶ�}��|s�nlܶ�;bK{.��;�e�T��H��~qr@���蓣G9^�ԑ�{%?�nIU���ɚw�@�9ėRjc�=���7�(8��	���ߟ����Q�/_�<R���U*���!鈃���9��08�))EJ������M��wyjk����C�;����Uzc���d�/Ď:�'�ԃU��%��Ż��4C����W�|��s�{m)�a�If��!�!i�����:����n�7$?���ʪ�LD@0��w������>p����
P�W睁Q@G|y���k
���'��.\�x�/$<��Wo�T[�ݿ�]D��̽���xP�Ql�,��LA���ǳ@���WW�23+$?������3�
&�W���!\12���N-�Ug��Э�~�j�c(��5})�A���
�l���>�i���g7�O� o1�];��u{p�Ӷ؀����!�[))\Ə�?O?e��I	�wNܯ{XX�8��u䏭���555�������BW.�sss�t���'�	W�$���HO�V��m� F�-Ӊ�,��BIq�~'���{$K02ޝ�L��.�C�=���� t�	������G�6��N�j��M�;��w����i�����*(0Nx��!�J����>^%�:U�f� �0��)o�j	�G
M'�ą����b��

��,�?MAޯ\m��]S|��,�E������ӿy��uH�~�d)��=��K�r�����f�>�������/g�	�����H%���|�u��K�~�/$4��Y����^��g��.�Ͽ�xE���P@{�A.��x}��[�Q:�?�P!����,Ŷ3v_]f$��C{��*�
˞Ĩ�H�r��� !�o�}Y4A~���IԤ�Pmt��d��$
9�����uʹ?.h����:Z�5j=�m�1;�٦x�0�#xPC���]�ӧcZóh��#�ƥ����޺g[n��w ���p ��xVj�"�������B3S�X�a��d��-�m�jK�Ox��c�,�ĝ��"�����.w�v�ĳgϾ�c��%��6)'���R��{$8��7��Ew��"|Ww<�d5��E�od�������A�s�)�Izjs�!sss_E���`���/�{�79� !����8�3�����J���ϛ��_�c�xy���xC/^�W�AW��ƍ��=��e.5�v��&�>�X62E(��g�sx�j�m���z@��۱jR �����J�/C��|?duq����(�n@�F\#�Û���ttW<j]Q:<�k��;�)�
p�&��[|'mq�n���(�E�Xֳ�'���%=M��nBd����p�]�z��fF�oh11�>}��0J����P�+�+а2���XE�@���ݴ���8XY����}@�6t�� ��3%���X�s{�ՇRR�e�U=�C���S�W���q.$u�gW�E�䈊e�j�;��^��	�=���4�|5/�!��D�䯭@���7O��/��Dv�l'>�e�)�|����Q=a��X���C���	 �x@߲ �M�T��e�������{��Q�p\�0<탙�TM`�����sT3�h��(��j0�y]�xHE����gM��,�e���L���zggg��8hj>�j��g�}r$��S7���'{J3���
@eH���$����!!!�ȗ~���TBKr�a�˄��!� �kE_P;�*�dU����G |8)�@�a,��������K?��Y�^\��a� /�"���~��fp7n@
�}p���~7���`�!"r���O	�f]�*����N9- ����H� *���n�n]���u��u�o����<�������_�&1L��߾b�Hƌ�~@�4���K۷H�ur�
's��<;[�e�*66�7t�,5L�R��Ax���K�4�~nz|e�����B*!
Iȍ����3w�81�J���u�uk���)z0>�"�/���86=hSo���C�KS���^�z	A�� 1�ՔHRS6�mB`D�SR�CR�p���m���a,�H�Z��QlGY�z�Jmk��4鯍@�!̎�����z��(N3|�2�-)x���#���o	\�OYK=����_-�����X;W.$/�̰����Ý�1O��5�=�	~U�꩝ʓA�O��A�Dh�t�B��`rx�c��q�'�]*'�2���톴��&nF5�,` po���/�?�7�	��ujN�Q(,.~�;�K
<$+�*vZ�J;�mX8R����̬��]+��"��w���R�7ggg?����;q�$u��� n�W<}�{�6�}���"6�_��ix.�y�F��n�ӎ
�M�%o�J���/	ȗ���PW�ܜ�\rĳ�O�mȫjv雙�? i��s�����o���n�u.�� ��=��<���'fN�*�]�2d��NR���Nʰj�.���&v�.ո���AR4 i॥��ٔ!���{����'	�OyW������������P(��������6��ze[sNc?my'D<?���B:��c`���o�㜨��~F�N�^�c�qű*gV���݊��]�s���e��|[�*���d�� X�<h��eBҪ�w��Kldd��T��"/�R1KxҦ@���:�O��_��Z�'P}�}��G�0��0��頩I�*ٚ��^me�v�]�t@R:$��o�J���G� Ωw&�Ъ��E� _ &px�:�������A�����-�l0���Ӱ�����p��9�!\���W�����"���nB�W]֕良�b����߱���TT /
-����*��á��Oe�>/ܸ��~m�#W'���Lj2��F�g�Л�	$N3�oڒR���@0�+�_�o@�g�$�A����r:b� �S���M]i�v��F�'*f%Fi��'ϸgF���ϣ���u��p��I⛙x1֢��
�B'i�8V]�.�>�Ox�1�*.����P���q&��3#�?|�K�2�1hj2�i���9�c]WRx~sZ�s'W���\1�f��Y�2�ǹ|�<_ꛗ|�Y�*���_{����Z��!�_�»�,U���'����B\i=�B��^3h�m�%0�f�8��{�ܓc?��z,,���밳�;�b���_�!s�L/%1��ꈹ<Jnf�.sYkw�(�!f�����:�7e㿸��	`P�ً�f\D �g��~H�v�=�=��&��&",?�����vD���R+l'ܔA���q�%E|����!�ް� �$k��6Ϋ��S��wn�2%��*((|� /�z����O��M~f�D���qB�ԛ8���&����Fr���B7F޵�?�6�p�����b%�C3u ���@��л���1؍6��t�@
Z�:����A~HA@mG������ ]SSSKdͬ��P r�����R�*'8��H�<�cH������/�,��Z�NP�4���=���p���y��[�K��E@Dd��Zm�xѶ�X=�N�v�ۀـ?�rR��G��Z�OO���/_��fй��J>4B^�^�y��);�Z�ց����T$�̓�lM8�ɤɧ�63���8 N�&	@?84T�r��I*��@�_�C���&�O��ߓ+;$Hg��YX�X�s-�]:N�(4�l�**WJ�x��6vs�H-�~�y� Z	xz���~u�����Ċ/�2���K�M�4�ۢ�bKkkH�
� )�|�$'c	�T�,�4ݤှ��R�:.�44�)�7{jg�������>*�#:Ǳ����Zƒ��G��U�2f5�3����e]iW	�Nx�@ ��<�8/֧w��@SC��T�8�;��	�J	2Ȋ5�#���{(���%�K��}|����_����A��G�~)V��H���ߙ%O�?�����t=N�>ks�Ǟ�������y"`�k1Vʘ�sI��=H�pr*Y�>���!v�x��T�����֪.vǀ���S����˯.\}O����N���.V�����v�<ħ��ɓ�;�|:J�!����
�����F�G��x�ڥ�ʊ�d	�	w���RRD�P�;`���]Dd-���'��)r 1��b��	XǄu[?�83���*GGǓ���k��D�:Y�'�����*ES�9��i�3��+��A�.��S�\$�����*l�	uN9�[����κ��gz�X^F�GE�^�����2;�J377W�ݸc��p���3Zg,:��B���$�C����3^�����͡���~�j��>���҃�Wc�\�N�{�+��i++��ǅ2o�y�9��(P}w� ��Lt��.����ҝ��u0���������HBl���W�޾{�X��F��4vb�-�-{�5����s<����#�����ܟ)�r���*�Ǭͼ'^�>j"��nx*뜑��7I&��=��)�>B�A3xy�-��Aå6�e�**. ]O���P,��4\��9�s������_#�4��ϭ[���O|�	 �/o���GFz��$�7�yg6~��R����/_r�3ɽ��v�V����545͈	��{VCMTx�J���e���93�*��Q^]��!�G	����OMYҸ�߼qi#��H�zOa��X �\\ʖ����'>�E�UN�hÑ��1�<�1y�xHfv|܀�]X9yd[8M�e�'E����T��h�(j�\�4�YXx� �=|��㳨��C&CIó��gΕ#��K�?Y!8�6���d�A����dN�p��HiC��3爕�k��pp��(�x���uf�𭸈�"].�>�46�JyN�24sGQI���u����^��>���%k��us-0�D��V����\��`4|�QF��L���DBC�C���ugq\�Ҋ�Ca`�l�`���UR����U��,,��Ͽ$�
�L�$"a�t>�}���Y�K�WA�q����Ѓ+��OX{�9))w�$��=��\|_VVfOAEUá��>�J����U�Ϝ���@�+�M4!����?��g_�HՑ���i�U�K�������X�U����Y�Qs�

� 8>����w�|�����Dt�xG1Ԕ��������胕*�ÿa�7�����ApwIi��X��49��C�I����� /��%�1����h$?�9YY�I����%�)�M��/w��\�p�e��)�T�����H�{�C,�T�&��t`���D�SW��<�1���� Rna�j=�LU��Q�Mϲ��Mg�ҒU�~��;;wq��>$�gr[�}��3�/B�2�w�g0R׮����;��>��[����xJ*Q�u����%%�[�ۗ����#� �I�P;�����K��)jK��p��bZ���H�{E�K�sss�8n�SXǹ��"��H��}����5�ү�u���Ӏ�~��t_��Q:�A���d�0T�^8� K�%v���Q����Ö��5{@X��D66�<��]��W� (XH5��FU��4���H׌6�9\�M�ޟ?�`�uk_���I��*��t�Z@�3��<p����mXa�X�]��R������J�$ ����
���^sY�B��wR�T;�:���6N�&_1s�ǟ���R�OsA���V�~��]�{��2%�qt||��S��{�j���
$�k����. ��Txh��Wl�l<=L�>-Fc���zo�猌��g���9�TI�w�F ���$���3��utt\�5m	�$����H����ee�̴*��QB +���{1�/�@h���.}��ɫ�5����=��o�RkkjD�=6�c9��b��"]]�wc<��llV���&���k.$�tı�D���T@I������+w�됶S;��ѡ%Ņ��=K�QOz�X� ���������l(����`>U�^����.7v�wŽn����t�!((����S�MM��cҼ0h[�|�F��7X�̽�#Y	J��)��ʚ��M���5��^2#L��̀ �>���l
8Ӫ:�fd]����;��@@�m4�qZ+�]^_��/��f����ˌ�5-����,���0P9Yo�mT[�M{Vb�Ȧ��j1��ͫRA��I���L5}�.�����H9XAV�Uц�Q�D� Wd���^����9�f�q�v���4�E\3ݾ���ߺ�1X�VQ�dϐC�U�h��%�'w��9���C:�V	�o�A��UK�ac�IQ�vՁ�4�Y
���A��փ��yyyw�ih���=w����Gl�cV�r㩯eךܖ��{���&���%jE>�C����%ĔP�[�E�Ϗ?Nd:;
���a����d7�õ�i����*��6����ni��Z}|ZP}]�.����u�G�m5������A�{�����ʌ�L���ƈ���}'�6*�8'�X�v(�+U6���}M#��k���ׯ/�!NO���fT�W��$��F��)'��zu�'�Gr���t��+�j:�����ې�n<�}���hϾ�D�):I�[�����]!��u[-�x���
l��V#<��3v֫>D�6�1�$�짫����X��W��]�j���߾OV��A}���y��{��v�o )^0���n�:;�E���H$���N0��7>�֗Mո\vf��8��W<Ǆc"
V�au@�b�.���&@R�H�aD,3��מ�\��!�����Ƭg�܇��5e��H���ꫵ���#:�ܑ_>�S���b����D�9�k�{g�!Û�N�R��	7(y�[����Ɨs�.?\���v�,;����nqrFu��X����p�ier˜b�^J	�:��Jҥ[Z(�a}˫�� p���ݶ�C8&r��)�:��y*��	���i���r�0���Ǐ:��`�M"*.1Ȇ��۾fz�3Ht����u~;I���1a\5���\���|�C"1��F����K�%���[]��}T�u[�,Dg�س&y2T���\x���g���-�W�U�DN01�I��g�Y���r��OՊ�������P�C�$����y/ @���.*��rD|���!h�n��y���l���[����ݽ�����;���9#C��tg��e�y�.WO;4_��{6H�'��A$��@�I٘��˗;���7�EH��K@V �76urqb;��N��ԥzV\��Ҝ�]]Q�i,Ւ�-�@'�U9��3�LI�T���'�Ɖ��$�u�k�MH;�10":�U�����멸q,xhE�����X���WP��raaA��|�J� ���/Y��g��Ǌ�!�����Q�BS����0s��p���T

��cRX�l�Jd�Zy5�� ������������-à1E:(����<D�����T���Nwh���� ��3ғ\�Mn_I���"���U���K3��lmo��+A�V�pLh��G3*�M�J�U��ˇ ��F�4��"�:�T-�}zz��bkw���lEe��;����5��\�j1���ڣ��0P7����vW���q�%���|�����""��7i�ۛ����5%�s�w�8,�I�����H]�$�='W�߷�̻��g����٫*))QH/5X8~�U\��X����d8�k��H���	 *��@��ǟs0W�b��[&�֙�ˮ�o�3Dpspx;�h{�	B�ֽ�w-e��f�UN����h�o�FAL\4��;(��{f%;r�����C��mmf�tAZ)��Y=}�v�؜k����;�ύ�>&���G��|��SXn;! ��+�J���Ўs欇N�QvFU�fmm�Y��������
S�����Z�������P��XO6�$�-%���ñ<f,��?�a��Vs����|0r(���@F�4L^�tl�"ᓰ�g�0�sk��H,�9�t�߅Ei��("J���d�2� �ڇ��4$�r��Y���%'g�����Fd΢C���g�ihP� '��s� 3q�W��pK|��H�P2��ҕ���M�@,��>��?�z����j��t����{�1Q���o�A� D5q�#��2�j%�6�Y�%}�ض���m����֋_&�@��CaV�����7o(��-,�999�,�֏{�Z����;������HWi���K�pU,%�1�N��������kccc�5E�~ܱ�cm%��{xCTPC-mmk�X��=�p�����I���g�Е����<<�� [/��D6)c3S�B�MA4� �<�9�y��c�c�^�r�Q�v���_����$�rh���;���>�^�^9�#un8;u�V*|�vqq��eY� ��(���^;��a��.y�9 d�e·F��"�������A�P�������n��q�=V׾��;�)=YxU��{ju�t�]瓺��"���
�+�\c8%�(�˟?7v|������v�<Z��|?>n��
�f�v<'�ٜt�3ǫ7YY��M���:���G`{B��u�q���~��S������
[CA�v&������c~�>�y��Pٯ�}���t��$�,���Ҵ`bxV˃��).jau�����o�*U/g�{�}RkziR�%��Z�ߵ�kI޿C>DGSc�deᣉ��Ov�s�*�����Uub�,��6,q[3���,�RY������wvD: :�Z6�^禨�,�)'�]�X�6([��=>8^���~:~ÿ�[OϺ������H��:��_�GȜC?�A� �@��
�!]���g�I�r�tg�[��'O�E'e_`脶�ۄ	���[^�H:�}�݄}c��uw�o�b��S5|��+�Q��Vo�ꏁD��pK���T�h���2hu{�ey�ޫwm���x����j�V5��>9y��u��ˌn���H�����vNN�7��I�H�ڈ�[d/���.^��zfn�0�;{V�$j�bw������7�U��y�p��&k�c�J-+;�P@�}$j&�������5r�Ɯ��;to��]��ƾ����O�O�ﮎ�J�_�IM5���A_'%|���_�ƅ�Я_�����;���L�ĪA�]�'��1�P`���,b<�̢������."�W��%�}�6�S_�V�|�p������Ssbu�����xؽ�@�ʟp��%ݱ|cnn^��6��>٭�=}z<����?,�|t�jٱ����j�?�:�M���\^����y��C_@�'9D�糸�gI�9�*��7An����,�TWw:��+o���N���c*�5�OB��A
	�b>Qa�ah816��$lb膤(��==�&��z���X[�Y)�\�K���5ܮ���G�O���oz��r���b({��)�N���w�:�*�o� ����U25M�MMN�r>����3̐I ����%$&&�����0���M�����Wi���i��ɉjjj�Z!l�p/K���c�b{ȣA;ʄ�z�`d<���$mU��\l��r]d�DK�Zńyk(�)���8��3����`h!H�(f���z�x�N	@�[.�U��'(�j�%?<�Lv����N�Y�I�A��p���bԲ9���$��scS�b��(*)�'�?���d+�O�oŽv嵵�3}IZ��Ӯcnif�|�C^�m���wZ����r>h�W󻃃��o<�t� ����M�&ې�S��-�Y);��ȆQʶ�L�o����vQ@�2�������\�U󫋇㹅ԗ���3M�í[ַ���{���B��~��Mn�$���f#��}}ʔpgV���A��;y7y �F���kZeK�^�ِ,N�®�@�}��L
�s�����d9������+������Q��덒b}��'n����__�d�77ݫO��=���g�6v���n�����@����CK|\1���?�tt��>�zo��#w<tR
n�q����!�w �>�Rs��ӛmW��������4yм�=�D0R-?+K�S��V	p�"ў=*�k�nݲ�I����n],���(&���ܛy1��drj�yN����������&�d���SNi�o�({l����v�N=+$b��|X6�SL$A����Q�:N��%����y�U����33 ���Su���@�t�ch܍�9��C ���2���΃���6])fܴ��0	>_�7N[�>Z�$V=�
D�S��m��G��J��G����N ��%�Tl��@�\�r[J�?�P��RK�����>��te ۩qz���ּ��2f����Y{�b).�k"��(v]E7�
���0q��[�v�?G|7��<"p)�o`�q[׽��Qi?YS�y2��n��/���T�jg�3B�+�~�QV����2�T1�U���1L���9�������/�1���zS���P&ι���T�l��i�߂�f�+2�=wV6�޲�8�.��,�w ]EE0�&�	I��݊<5����D�����c���\���5�+T�{Ǿ;;T(�DhI�I���4�|��ԁ�Ӣ�4�������'���;��]�k�Ս����'�n���1bj<�\���iy��~zca�&Ӎh �č����ߎS��	�+�+'�rp���O.|��gY�(���`C=��s\�k�?�
�?�))(��<�q����z$~�ur0�ȥ���\��+n�׹wϛ�ٳn��=�o[�־�������� N/chX�$H����.��F\��z/��}�5'Q�G��d�;��}�LKMmQE�mu;�=��[!��Z�V�� m�/���m�B�����^�$:����I��J�?Ⱥj�6^>�a�7.���ϯ�Z���=U��D�!~�3���b.�/x���[�V���F�n0:��0D�,�hgW���j�;���X��a�w���I�:�E�*eͣf�bo��>�J�%��}������w���J� �m�=6���훉���0��g��.d��T�����s�?L���0�����<���Ŗ=�7P(w�W���/��KՂ��\�e��ݽ���4T��j'�Ơ���q���|ㆇ�zq�:��<�f��T��&j�-��Q%οTy�6�&�O��ȢA������h�MZ��Yz����q��m�DT �w���[ٻ�N�g9d�)��8���B�r�O�!����OH��[�����LI��I�㡛8��/b�O]mllw<�<@ -*��7'U�32��Oq�l��`ee��^*�kz�c=�e�+iީ�Eƚ4by`^�#��k� *�-��`���� *�KV��]�)�??Z���A[)���P�i�y��P�*��v�Z~b�x ����~��}u�����\?.h��˪I�w]o������/&��/*��+�R�ſdGK��۳��XN�Ǵ�<�fef^L�m��0[�sj�=�L�є��Ɔ�8�l�4��?T�dEe8�\Ÿ)E�����숫���Y���J࿾�d�h�%��Xvv% ��ߣԨ()J�P�ǝ��˄�.K�
**��t����|��!T����+jX�׷!����H����4��ݟ���56��[�<oԽ���Hr59�Y��%�����,��[5�'���~s!�_c Ԍ����Wķ�ݧ������v���3�=�VG7A�<�O*�"�P��˄��ElÞ�n�(�i��RU�s�����[�U�m��7���H�"��J7�H���
�)��D����E��"ҋ�Xt�;o���s����p�}6s�{�_�9���N5��RNN����V�u%b�t�D{��������+�wo�����[b�P� �?���vV����������Z{6~�~ט��#8 8�g��qĺ�~`q�ܢ"�g{��%�Ƅ���@�8�]z�U�Sj��cj�<q
T�Fg�T���'8O��i�ސ��soB"��Al~�L���m����YX?$;D,z��u{���ڹHm�Ŗ��V[���+�Nrc���t�3K�BԱI1���ߢ�'1U	���h�m!x�C�EqC-.��}v�s�nھG��>��~	�i��Jж`�s�?��Niə�+�6Q��B`oﯬ��JJJnh1	�G�A����[����'L����Q@f��F֬Q�g�?Mr�Gp���酹f��k����L����S�iFm�ֿc�����@��(*���{��!UM����pP3���I�n���p�^+v5��))�1����4��d���ڼ�c�]�������DB,�>�{ha��;?���
�5�T�>^i���#�E�WL���Bv�\�p��|v���S���6;ZI[�c��V��ޞ';{�LP���^�s�888����H�/�����Y[m�k�C���`bh���D ��X���n���t�.����1��1�<N�2����zn~�|��%�����N@�F��˟unڸ�䮨^�s����h���p�v����'�^G��EE�D������.U�DM߫7���w*�5⻽��пG�0�i�O���r��il���~����q�Ѻ:�9>N$9>��	��`W���U���4(��w�w.�-�d'G��4�h:Z�̴?m��/�>�J1�b׽y�w/7i����k���P�m�|��]~�Ŧ��z�i�y�9�o ,bh���gA?�o|��T���|��.��U�|"p[�`R�Q��(5zG���ualbB|�mnaǴׅ'��8�hw1b��h����o:NcF�Nu�G[�EY/��/�E�\Z�3����
5������<}����7#�9�����x�^�4��@֕�����J�9tF��6��L���'$P��P�f�}wyk�=�>��E�K�0<ަ��	ăs���Ǚf����<�?rg�+| ��~b�쫴�8�B��S9ʀ���ʲ����	x�M�W�\�*J]����o��N.6R�m��[�`�k[�O����!`G���k�mx�X��'��=��>��o����Ɓ; ��[�n5	(X_0@��[ p>�_G|U����e��i:����;�X4�b�cr��8|Z9L k⾇����o��L7n����֦
�{î2y�-H�O`O5>GGs���j~z�	�������צ�Ո������9Q\���̗�����w+�p<0 S���;�.��l�b�[�6����"uپ=W�+�{��@�lE�%:�Q�|g=W���@����x3B^[�����3d��^��6��\��p9��auM����M5�Cy��ņ7.��:m�"��ߍ���_���﹚�Agk��8��Wu��57�^簢���Ȼx��t�������b|l�n4��#`$���Ş�[SI���Y5���pkn��¢l}����s/y%q�s����P8]>;/ �#�-,()��<L�~ἧ;; �}��T8Z�)�����ڤ�f�޵|f쨌���`�^ˮL�0�p��z�����{U�ܪ�E������p�������f�wtr4�Z;O$��T�B�X-��� b~��$ٓ������������r�,��FQ���Bx�G��ǎ�����9X�3X|1�U b�i}Z�d��+i1�ϳW����u�Y�Ro�I�2������e������aJ�>�5"�;���4���~"�p���M��%tT�Ց<�##C>��_�w�	�W�/j������A5�@���<6�<^����6O��Y�ׯ_I���!�$�+��LL��תYX4�>�������փ$�l��,9y�`�n�����=	�64��$$�rr�k�u��ZԖӍ�@݆���1SD�P(�iu 2�D;���q��R!�O��KDT��R����o�w��
V�|o� 1K���WJ��o�L5�ݼĒB�d�_�Rz R����5X��|�2'%e����Ȝ{���e�k�J"��U��&r����:��u�#���Ы�v5����:������[V�{�

9E�K}ꀓ:�\��Xܛ,�?nH��Z=�Іe>��:�T�����w�2�֓_	JU��ϋ'�i\�I&�5�><<��>� N�m�"�j;(|
>�8�*%�����[�w�H����U/|��X-���;F��@ Bv������������#��XX����c��N�,��ǽŅ�N�5��<�ښ�^J �����{�V׺��I6�D�$/t�^_���i?h�8㙎Y��q�~Bu�O �5�ݬ��PU}2��R�l��-�����T"/ v�/%؇�����y��zʭ��yc�2>~���c�+�/K�[�����ccc���l2� �ƗH#&��Ю.y �H7OΒ���@�: ��I�a�VPХ���礨��o@o1RD�Q��i�+�sQ�L;�\m���4��4�6&�8ސ�s�ڎ���i_���wp?��a����O���;E+�{.�571��wC��6���~�1�f���O��n^��� U��<���e1ܥ���y��3��w�נ���Kݑ·n;�URpy$�3�G�w�������Ⲹ,P�u� �Ng�D@mFf�Z�F�Tpn�޷���c�������w��Ց��I�P���[�ѻ.A�0�2z]�sSS4��c�&?3d".��,
8�]ꪢҠ�C�=`W�U?U���g�#�x�/?GL�x�o/t.,��cB�"Jx�&;�u�E�ؔ���P�ӿ��tMf�O������b�X���m�]�(U�tu��eH��h��:3I�e]OO�d&2�a$�o������*���b�H������o��LUW�����#���ቺ���K�)kQ�$t���0�ZEj�W逋�����QW� �}������T��~�fy�<���	�=\�"����=�jk����c��z�g�B/��� �
	A�<�_�ö�+=016V����3��U-x�|��S����Ӟrc����^y���6!���Ҧ��:1�a캵\���uȨ�֘x�gn��K����]w*JJ���C�ߦ���nQi�f��B�1t]N���/J��^Mv�{
7_���Q�[��^�e�����՟`��080���
�ݰ�)���r��kOM��&�{Fo�h�~'�g��_�8�H������*�+�x��}���E���&yJC�}@	?�dVs��>n���w���f�?�t�����w��&x:@����6F%u���3e#�UWWCʹf�%�������jg�[������\�vU
q�~��@F^ޣ|J���Aډ{�p�=�i}|vkk˾����x��)%%�v�5�<՟_r�U�V��#�$��}�R"w�ǣ�r̤=�>�	�	�Z�.o�%�C��6iN� жrQ��<VTh���#��(�ϥ��m��=��/J�BmQ�
%��X����OO��.���Ž*x_�yT>�?�.�͑��񲞪?���Kp����~1R�}���cӪ��PVF��=1.r��0�H��i������څZ��^�[Q�'hCLd@�ye�7����� %E���KÃN� �=~��w�!>J�3Iƃ�p�/
��Gf�7��BȨ<��8�h�-d�y?��*�f���(��b���Q���moq��ZΏ$�����X�ڰ� A��x�{��)#�I��.�]���l����e ��Z;D�/tD��l,�}�4�g3%T��#����Y'gV=� ���@B�� ~4�Z\��~I������������X���!�.���r���T������HL����	&������S۷o�*�ߍ��x�6��; �c�HI���ӿ�$
����(�ߋ󘮝��~���]�S嫖K���`ېK��j�5���?��HHH��
=���h�D-��1u��4�S/5hcoll�גu�\�����E.N�k��'2����A��ɔ�A�Ha�52��A���$�͜�Պ��h�>�G ��xo���zv�����4��ӧ�%�<�������7o�=<<�a s��4�Z�=rw����0����yk� "���:g��w�u�����R�����5����"j=�_��@8k_.��jW�}����70�VL�����>|��نý{��{�5�U����@͕$ֽԂ~(�E�6�[�T��@�W]1S�j-�͆�"O�i�9���s�B����V��
z�_�8�]MF�Q� ����ӿkU�~W�i�H�����Tgg><�*�P��jL���ڵk]��킘h:��7�B��P��uʙ�p!f����`�	�qޘ}��L����\�ti��%
����	ʏ� \�0�����ڿ����+���oBOBoK�ef��\����ѹ�t�fj��e��Г, ���Ƿ� �W�qdW3"؅��6{W��(p���Pʶ���[���ٞ���V`��́i��%z�Z�,�_��ʦ ��̬��98��6,�q�I��s_����.H���;��}����%;�Q�t||�����z<z?2w[5�}�v ۢO"���L��x��x�����1�C}�	깢� j�-�w�M���N�5�^"�F}�G�6A������G���C+�-�_B]�j���[�}�ԫ�C��ÉvG���k���T���O�W�y�V���̾���9�il�ŏ��ȈO%�� �O7��`3W�U(�k8>D ��dq"4�Zs`�Ê���'�@��v���AK���a�FS���|s9Mg�6e��w4kr!�9�D�t��9��~`0�f��V�� �!��*�Z4n	���C�Ѱ�"�;��/X�\���Mu�N�h� ��eu SN���lBJJ�`
(�l�y�����z��p�d�Ku���c�����w�{Ě����5�)�-O����<y����gH���l c�o9L��M�`Tc�3��K�ڄھw6S��F/%��O���fYy�0V��}�r$C2��� sIjg�7�X�P�'I����W	�xb�ҟ�B��b��K{�����[(Hɮs�vN��uY�@�ך͆����8Ե4Y�Q�k�����|�}��*�n�r��V���NS��n�111���� ��)�.�*��lT�YqMk�?%��oj<<v{�:�V3w)��S���	֍�29�L��w�ļ��� ��`�����
�)61�Ŏw��mmK�]p/	���EO�UV,�#N��p9ً�3�C�a'oΖ���d��� J��<.����H��sH=55��J9z�ϻGR��̽&�̰
|xW�JG[��p���qX����)t.���3��yQ�o4����#JhΥ&k�2��?M�3^t���ꃔ���0�Y�uu��\\�B�=��S�=�g WC3�;���y˿v��DX��N��a�2�IK�� �|�=���R=�d��Ԏ�g�� �nlzcf�>��:��~�q���}�F1���&4t�����'��t�lM N�0��m�� ��}�Q��c:%�c��&ɞ��se0[���[�"�>��I��yG���.I�O�P>` ��Xք����߿/��:���Ia���l2M���l�%U@����ȄkJ�+T�@�tma�و S'�Ռ�4@�'5�7�h��o�NU�z�P���D4k���1==�zuu�?=�kf%�!ͳ�}���Wa�][Y/`�#��޳��x�.vu����u��-����]�3���q��:�ȅ��s�XѦ"�P� ��A�e ����i��B[+�
ҡk})������i�ҔB@M?����/b6�jO����?�D��u�P��
i� �4��]�-ղV��@�] E��O�'��K9�E�f�fb�� ����{���8�r�G�Hv]��404����u�����~sW��>����=mmy񶑟}9�/���k���J�"���Ƃ����	=�H�؎�h����?UK��'�|j��$���A1`��RO� �]���H�13��>����Tm���)�s�=lQ����8�	���Ϫ&�wr സ����.�/������ ��h�7�
�5�y$�'�������Y����I�Y5�������G�D&�\��%���bX ���cRJeq�yˌ���<�8��'Y
����O w�B�����a```���.	�������F�3���D��u.U�fj'�^]�%���짃�r-��������P{�E�j+���� �	���F�:����G��bo�����kfA�սϪW?�8�7�U�OL6�����4z���go�Շ�ÃӮ����Y�-,p3sr�W�kR���� g��ɮ�8*�m��j�c��g ��d��"Ջ��l�
08�?��u���^�7���GjUcOP�������e���w�1�}���2_ݲ`�E��6r9p����җ�6w� rʚ��s�9���C���Qxl��UL��e��Uj�� d��N����H3PC�Md��6�����o�sJ�F���[�=�:��qXa1�xzz�aZ�b5+�=Yg��Tnn��mF�E�U�o���|jV/�^W�~�?��E���Ui.��-̾�@`j~[[w��T�yRҴ�P�@���'��_�7n}*))9dy���㲵�_�cǉJ��<b�*��E��V��6
	|��?�%�E��K�� Zc���������*�j}��
��4w��~/��C9��QG�2�B���k"mS��ɡg�\+i}�z��D5���%��B���- ��c5��H)]�j�g��W4H��"@2jI����wEkjj�~��E�j888Xppg���a����9Y}"����u�9���)1�)�(��J. ����nIJN���8�W휲��g�0e���\��[����逽+�G��9�ѭwy!�<m̥�b=����]W�̣���)@�*��5ww�r*Tbf�r�Gf�E�+��`�K}��$z����!�����I��A����J�Dz\���N���C���f�fW�Q�%<�e=�
�j����l6�`��ib�m�3�=�j���{��-�Ϫ��R?���J���y�}ȁF{GԤ'�d^d�b��������$�{�r���q����6�j��9J�(�j��s3Bo�� ���5�1��k�ݙڔ�·x,C�v�䀡�B�a�j}<�<�2.4���R����h)���ֽ�`�]	d.#�Ц���C����שׁ��R�3n5\���!M�2YW-q��.��S�a<��t��������s�B�.v�X}��?���@~'�QTl���\M�cMrLT��9ȩ^<ex*����s%z�L��S~�Б1�[��
�|m�����:��*����o�Y2X>~��Q�����rc0����{	�1�h��}�A��u��7�:�ǔUT�g(��	H���g6^�D� J�G��O���bBN���#yd!�@�s.I')&�,xZO��.��c�q��P�p͖�I��'�`b�R�qZ@�*^"�2u򔗖�'<��?ߟ�,Di�o	*e���x@>IL#th��������O��t�g�_t�L7�i�v�c�����ur�mr����V
�C(�|(��C�������5	|oğق�ʡ�:�We�o%����8�g��M�gc�K���t��q	��n���E�##��K� 70q��~w�D���
��_�:���I�A�K�Ή[�|%��5q{�rD�^v�i��P�X/<&���ʯ��/oێ����<�CMTZ����<��F�O%� ?�E�
�_�w��	���Y7J�UVr�ݝ�E������G2��ӽ�l$`uC}����V������q@�U�X@Y������i7QF<���刁�adcu���쾯T��s��mR��@"�Q��\�J� `1�����I؝/�,'��)�ݸBDDL�S:0�&r�X��߇�9�����^���vF����|��P�UPR��l5ܨ�"u)υw�8�C�W��E8�n�'�?�*ͨw��3�}6��X]���&A������VՓ��C�Γ��{�#�ZF��SJ��'l2�i�zA6�WQ5?�ZeH�3�x^Bd䞲��8�81���=�]]��@�)lK�͸��ډ~s�c�\��rr���5Ԏ�7e�%��.�����Ě'ۨ��e�su�3��4ɳ������3�KW��BC�dc����_��OH@H��Ӝ�K:��|�)/���oӨ)����j6-��3�U%[�l������Rf�^��9^��&��3b�TS=#�"ǂ����7bN�6-�5�%'(E��
�mG~�b�E!K�V�
i����#��>�F��?��.��W�$���qW����?��>s�����W�	�%��p�=Bo����Dâ���w����L��T+A����mK�^���������}�WZ��FC��c^|�Ϛ>����9�7� 	�|�u�G!|��͛+����΄7�Gl�ޡ0����Ƈ��,��gkκ�@�B�M�7J"$�5�}g}����D���^�sz(�bT�����ӏ7�i�D���c�O�u���;Q�Y1�US��L�4���,3��� �xLi��~ՙ�~]������"rotd"7&�H�ݱr�^�a�}�U�Fa6��0Gf��v :Y[��<��Z�߁U�]��c��%�Sc�zP�.9���]u]���h*?���ћ�o_��
,����ˣ�e��ׯ_�_`Q��S!mg}�l332p�����N�������~���/�I�<$g�h\Nk���T���u�ݩ��֚��h)<� 
U��| \C�|����M[�*�ص�J����d$�����e�/�����[���e&����ͽICI�q��%?s�� �7i��^��'l�U	���lm��L6x�&	�݊�ӵ��df ϕ���,�E08��l� ��$l0[)�7��*&&&��z�t�o�_:ԗ*Az�#Soѳԯ$�O3����xC_���t�ٸ�*�iS�u���s��g���op~S��p�x�=+i�������$���ԍ@R�����"�b=6���P8����B�jg��n+�?Q^g::۹���5���m���g��� �����'�β�p�ƍ���,��k `Zj��YX,*��7��yiIzgԲoNMM)�͋;��j�=���Q)�+3��8�������o~32�~�xܝ ��x�-Gjǡ^Cg"..���N��fj;�ҕ�B��G[*Y�cw%ợ��4�݃�Q�k\BB�zC���u{ �$d��:P?��9ے8��,���h{��`�R5��E�C�W�9#E
��K�{�@^O9��%���@�c>� ���=F����Vx3�Ց4I����t&�ŀRDE�C)%
1��#m�L�_�t��<}�3{vRPP� �D���sg�����URJJ#<1,0���8�jn���X��Hܳ�#��D�ŋ���C\;v�����W@�֥Nӎy���Q������frݒzY��V���ћM C, q���-�]B����<x�`s�˗/��ܿ��� ��;���G�A����I��f��A�`��F�jk*�%�}l	��bKP-K_���S�� � 4���f_��yR��N5�.�a}<RR���4X�� �a6��\j �m�B;ajїⓋ.�qn�.��d���Wwi��P�[��m�DQ�q��45;�ȥ��2��r�3?x={�,ñ:|�"ߒ���n�<{��"�qɾP�<��i�l����SbVN���tV�eRI���&�;��Fgϵ��ӥLD��_��m���e�ٽ4��P��è�(��Q���X�z��9A~U��R�p���FX�gl�x���oO_�k�S���z}���ȧ�ugr�/oCݏ���Uc�1U<R*�kxi���=q�����؋�Fܨ�&�sU�B��
u����N斊�v���S�����i@v��˺�����Q8�ǃ����66����q�[%��	,��ٳ߻�����}|Q >eIr��������������g�
��3����eE�ˆ��҇��
.�8�Pk�����Tq��� ��h�P����/�Ƈԇ\�)XɎ}�|Rbb޽��S����� 0"[��\,6M	?����� .���ˠw��e��JD��Ey��v���ׅ�/��#�՞�R=�2˱G�D����v�������� րm�6?߳���T�c���<?;Q��ΏZ��TZZ_g�h<LC�0K��n������5-�_0��oD�-t�F��b\.Z?=�YTO>��S��"ђs�nչ����x�{������}��\�px��a(�����F��[��he��tn�ɺ����IӁ�7t����4'+���^�P�
��]Z>[���5nN���L�Q'�=4l�(�Y"�re�R+�Qc�[}5��'a�6���C ���멻����1��Ǟk���<49ׇ(,	��
�,%-��_�Ezxz�k��l���'g�A��y��K|��>;���4�B,�hi�x��r-��O����$�o��M0����E.)�_�3D�a�胼����C:�/��:.���E�B�}��*�f���'L��m�dQGOZ~��p�������S�)��A�M��|�s��V��>W_�H��E�+�B"�s���c_�Ȯx��ޞ}�zgƚ����Z�M�K����qϸh+h�~��8����S�>|T��@��ӧ����q"III~�A�Æ�j��)G.���'�)6�#a�r�L\�ח�'�<zۖŪ��ˏ����"n�^,�J�V�O>�uq2���+J	�����<����̹}���\�Ƽ���<������g��&//���B�Z��# ��
�1e@p�8X���>X�]�^Kq�Ҋ3�]⫼Sב4=���m>��/�Qt����gr�cb�3~Z�\Ib[�i���C0?�m��i�c�糶DW�E{�͘� �:����n��p��EON�?�\���7����
ߺ���d�ި+� "jf�3woj�(y���w��p�8Z�Ȑ!&C�K.Gd}AQ�^��ױH���Vիw)�����H�*��>�m�;m�*�2���_�h+��e���Y��R�x,��'Rc�u�0g�7w�6��c6@\F�e����Hy������ơ\�>��@ہ�#Kn����u�+�o �_���QwY٧��4��kW��$�r@)��iEtDN7%��k�l�vZ��&��ݽ_�v�Iv��V�Qg(� PW���vS�[�s�?	/�"��]�v,4������m�)ܪ�[(��{Ǵ�~ Ƥ�!ԣ�a!k!.a���!>���|4 ?�ګLzi\/�)��.'򑆺� �R�ď�.2���^wg��&��?�a����w��m���ncKKl��Fo���n~we��vV<b�E-�3d����p�u|x�[Ql����ӊ0��y�2��Gu��D���9�pj�g���u���c����8��s�&��f���ܮG�B<��[!�$-*���׎E,4��\�d�cď��� ,!��ɽX���g��J}}=�ڬ�f�'��߇/ȇ�h:66���{5�cgQQQ�P��gO���S�@3��8߀Fn��SMLL̞�-�e�������g!/.)�]��d�f��Ԃ�k��	�[�i�A�v��H:��%V;w�5��WFھ��p�|�X]��)\�{(l��(fX�惐<�?*m�E8o��@����걂�E�y���o-@~B�u,����vm���^��N�Wɒ{�8^�^K�i�6گ��Wy����cŢ^p:��z�>^	����~��A\��a�n]��|�������Ge�]�ݯV<o�(�N6�"��fͲ��<�~��~�Ϲ��k��3�� �w���Cw�ܙ�YJ�H���+�)�ztQދ�>2�@��(x�2��{����vt���Wq�t�6�HҽLx��s�n�6#R�d�x�v�0AB`Fu��X�a@�!-������J�99��i�����_u�k����|�*�9�e��~�1������y�콘(]���,|ސw��~{^��ZIF�jgv2��ܞ��kaa��� e��U��lr������a��V�����ۙO;O:F	�F�l���{����&zDf��P&0����@wl[.*`���/YJ!�c���H}��4��>b��uΩ�MN<R�I�}� ~r�ξx��[`n{,Ӵ�,$�M�6!�|x0���!�b��L���/Y ���#`��{c@��ނЩ,SN�x-wa���21��H��mѿa�-<<.c	��mSv�H�2���ӧ�4��x�8�(1J,�O�mcG�K#��"��� ��ͤ+�bX�����R���:'���G��J����xw�VX&��+������bD�ˌ������
�f_z�� q�mxF�!��������y����Y���Q���R{��^��\Q0Zj�	�d�g�Ǌ�[Z�㺍Ɠ�@1���{��x`p�Ծ)^�,�����~�/E�o������D�O%G��p}؋����.�@����N7z����[�j�2Y6�ܟn��₄�2�������.HCGF�2~����8�����Z	 PZ,� ���^k��P^�8Y�r���pw3��E�'�k�pH�����#�����s�F�`�z!,�S�ɪ�-. P"��V˿TE����T�D�����rls ?����2����H��3�E�<��t}���tI����ŘU�o���cg+�R*�Q�ɷ���%�ZkV['�![ʯ�~� �z�K?Q���̲c��q�u������Ƴ�07�U��M\v���6�0,��Hb{�[�LI���Q�c�H�)���=��J���T�ns[^^6���
�嗮9�Q���B����,ݞ	��UP��w�P���7c]�(�}t�޵<#3"��!����V�����`���ȃ1f���E�,��$aw��^D����T��9�`����%�\e����k͉�T�`P��4�0�,ݙ	�������l�#��o�l>��@���OrS�@#�13^����?N>|���9��X���e�f}��r>+�:p1�hC�_Xo��\�#�-|�ԪP' �x}֓�O��h''$� ך�����P~���T���!1�����B#4z��qcJ7�M�X$�	�Ҭ?���ޣ���	�f2Aꦢki���Ց��'���ķ	�� ��W��M��d���>>>��;�?����8|0R�E`f!P��${r�L�V%nm��]��B'�迿�ܼ��c���Bŧ�����<Kaa]�����N�_��!|º�{����!x<�����|�+�,��@��,fm�����ȧScg��]�����=7� h��5�-7&���v ��\�:'+�!�����j�Q��̕-����m��AMMM-gj�z���X�Z���9 ��y�.fce��GG�([��[L]\6��6g��T�A���A��c*le�%�#_-Qe]�5I#�1`��싾'����A��!�@�%�40�	�s�D�;��8i�1 [&l�ȌWN~n˩T�|�;vǻf��g\\&��3��=��	�/��+*�v�ū�h���\��~�&� 2jj�*���!��
�p��l�6�.+,Fz
�;}F�Q�,t���?�@���-w��J����o����N�X���~���غ��D���+�?��4O��̗h���i] BЍC9�*N�r�z��@(+�P{k�oζ��V<�NJJ_#��L_P�Tš���s�k�v�zy��Cp�\�w��L�H硤Ue�S$��K׀l�愣-!�����q3��S�Z��Z5�o���ύ7Y���\I()M3����sv~J�R2�������1��,pq+����|��{��4P�d#��w�60c-� ������+$�:X�'gV}�6)�K{��ˎ���&��������+++�8!���p�+ �%��Ь��Ek *�Z�l�%{�P��'?~ �2����G��
��ԭ�)�զ����Ȁ�P}����E���hE,�c���*�_��bIѝ���[�KX��ؒ�߸��Ċ�>��w���~���7�o.�ό��\�FVC�����X�oa:L��;!Wn�t��a6o��I7u��v+}���֓B�AA��|q���(v]� �h��r ɐ��/R�=�&���E�� ���E�DO7߂H�~�\Mbqǉ~7��F؜���tm�T��lë��Xt��9�Mv�#��ŷ��l0[I�a��t�d�q���ԍ�ѿ��w7nH��.����o�uq�S�F��/�o �/ ��Il�;fFZ8.�T��=�<,�,7��{��pE�0Q��B��8^v��B֫�t�#�T(��9����P39�fY+������B64�'�;��#_h[\�+����д?M9S�|>�O��� B�/^�D�k>��A�S|V�tA��ʀ|�X(�%��Z^U���g��'�m#���'
������z|84��l_��"5�#j�>�ۀ�; G��9� �B9K����>�h�������Z���n�ݖݡ��i}�l��X��>�][39�4�M�r�)�G�c; ��S!�v�I@���@�6��8|�@雛�����А�{չl��̘}a��F��ݙZ]�/n�a��>��*��*���Qwo�RG4�U�*K�"5di~9(�����f����D1���q� �w�=�(T.��k�X�1�pa�J�0q���*1��.7����#�F�6�|c��K��{Un¥f�I�]X�=�2�����OQ7XCBV�+r�յ�Ͱj��	�J�N��62�������8w��6j�N��"�,�˗�;�$$$��� �l	���d��̬s�q�↰[�<�1�8��[B�����)B�.q�2�Ǒ�`� N�N���r{�8neK�U� mYYY�
>>kv���0��f������,�pA���\֊��(�~��It���Ԩ-�u\��#���Q���chN���h�����v�5٘_U㻍"�|��uu*ھ}�{�yg��::,l�C���rk��@Iݥi,�=�X����֧Ih��3L��(yX��S@����π҂i�ZO��`�G��"�h�`������f�J��g�@��D���3�Ix�/Z8��$�D�$��$��� .���+� m�4؍��e��}[����=l�;�и��¸L9U �����^8ߘBb=�~~|�gZ�����P�	��x�ɖ#��<+G��LMM�&��`�4�Uw0���?Pi$��+t.���?75]p�r����Y�/==h6+Q��gU��(���}��y��׫��}����cK��p��<��Dg�E����]G��Y��u3��5�y�Mk�jS^i�M@����L���J*��������5��,m�ՙ�)�_��ꑹ�hN�qq̔�:0�+,O��B3߂o����&�L� ��xt�P������	���Z��$�r���Q�s�����p��1���Z���T�����UO7G��[h$�mʚ�o�X���4.JAb#.�������ޛ����#�Kgf%��%��h�S����
��ɰ;��DD�+�<�Y��=�M͜Zf.��^c�od����^�=oG����1��:�9^-�|OBHl>��4���hi1��t���ԟG�k�N���	��Y��a��X�c��M�����|�����r�·��נ1�NE�� ��e�7h��x\����xD �F�NV�����8�n̤wނ�L}}t�*�4�F�Md	66vLs�����xن�(:�|�f�H��a���F<��@��l������I��ȩ�r�e��/v��*%#�sQNV0Xa@u9�If��Xձv}�R�������~(_�7Yrw���J�W�������~;���L`H{g���r��<4��3Aۿ�?�ʹ{Gw��1�`�ӓs����Z�t�����K�5��،6�Gh C���/�����D���_cc�b�x6Q��#Z@��nz_���p���;���t�l�2J���}���͞+��Ċz5j��@N[��J��^6��Ç=�5K^�@�^@�D��8^!��ٝn�"�w�'���&'�0�����A�w��lg}�j`�ʒ��|�P�b�3�#��h]��޹j{�����J+ҟ7|����6��	�y,���zr��6���̢��乯Y���^Ⴤ�&������q0^�����v'G��7��H�?I��ʯύ�����Iܣ��&c�ٿj�����W/�i�$��`#�V���6�u*,���~��6�2���X_�� ���ɓ'|?{E/��4ˍ?�5+3I@��U4V��3�s�����W�Ui�r\f�qٜ��'����[��ժ�S9�?�u���ivL}�C#��B�F�9�o�do���
yε�kЊ�
hb ��\~����R��h���K,/�KA��"��Ҁ�T�-~��]���'l����J�ͫ��`��`y���{���������&}����� ���Ԑ��U;g������]�#�x�0���~��d�p�ʝ��v�)�|h -"�C�����<r~>7x����I)鳒��IK�lc�Z)$K�� u#�B��G��Q4�{;I�����7����! ] ?Tb:$~­��2��Օ���0�WXj��ǇfC�UU?�k%�.�w�^>;��������rg�D �?��U�2:8�
�r2�~K��W��Mz��]~����Y�;a641j����쇢�@N���4�|{6��C1G�T$j�Ү�4���i:�jn j�h[r����V\�Q�S��:�IOLh�!���Z��T�u�6�$_�Gg� ��\q�J����ߗ�bƇf���,)8!�YY�X;#b�-��>cz�ت��B�y] � �c�%{g���xxxo��������}�]&�K����fT���xڀ�u�Te�/t�TӞ��/��$2ܿ/C���� ��l4/�~���
^�«�S�ګ*���5������V�������ω���g��@�'����˪� "��}������I}JJ
X��?�F/�A��q;�	%��Q#b�>����+�oAH��P���Px
��;&T�ϟ�7D<���+��l�>�|�ڨc���:�T����{��2���b;,���=�M@'�s߭������,�j��z�U�$��05פֿDG�� MІ������L�`�>�t�x����20e{@�I%���Qw�������o�HD���D�:�{��osr���r�������.��7�pKd�
\��Dr��$�fGh�4�u������$b{4�};��Mޮ��4.J�o���@&τo�ϟ�e���[�>2��u�П}
����Sc�	}��r|�����~������=�|��ȼ`���k�Qg�� �ԅt����Ǜ���pOh�^k�i2�YW�hv9\�f����w��Pgm|L�ݨV�[ﲱ��i"��c�U�u�]�RQ�H�T.Y��!�I��`#��r�\f��M޿�?�������<��s��<��s.�݅��H�'�3`w��RVS݋�g���G3��?����Ԙ1����^f���,$>m��X�L'q���.o�z���I���9�B P)��,�!�'+=Nkl�����ᮜcg�g[R9���w��0&�Yq����)D��4��+&���S��F6R�݈"*9��՞���u�ϨOҬ:m<�Uat�͝����[)����Tz�]Nx�E�`L��ŋ�(Kr�gcL���=�k���_�����C*�


���p�jU���ׅiT��Ġ�>�w�ĨClZ�[�{������8�Z/%ž^w��U��+9=-8��W-NBE�5%��4k���'��I�K5�8�7X�b�-V��,�P(�3t��`D/�C����"���c�a������)����}����}.W!�_X�(���'�y���;>ypxA�1P��8�e�螻v�e�k��.����YAaX��\���P�RΗU}��J��f�JK/2�P��d���!F�[��yo�ԟ�P"R��ԓ����X����wW��:���ics�������޼�|VT��}|a=����U������H�iݓ�T�5��ɂ�)�����TN��U1p�5�w���S���yj>5����c�I�}�F����%|a�
�sk��=���Ί�*+Q�d2mP��K�o���P6Pijҹ�m~��p�0�I521�>���](s׾ ��#
l�.tϓ4��c�x&���[���FZ�}�?d�;ccg��1�%~GwB>���ul�
�+��v:M���4}ۀ���������]��"��^�v�[3K���@
{(���*cM6���%$��5�j�Jɂ����"�QVV`��a9b�8z�6�ĕ��/[cDZA	�(��\�O�xɈ!���� �y�s�א��C���
�)̰����Og�Ko�ߒwvvF�h�L��f\ee���'�f���$����>�q���X����6� o�������e�2�bbSJo.W�^Ք��a������&�����n"X2��H7�ۈ��7�����"�v>$�c^��`���	Ru �	���?�D���@2R��mw�Ljӣ�6Nq�0������Up	��u>4���d�����O~�"<ڇ�a��x���[KW׌"UUj\tL�^fyh�&C򒜉���l5г$�"3l&ޚL9�|||�<�ϻ"_�lmED&E�;��KD��/�� ��]��{�]�ڬ�l�׿b�O�T����(IZZz��W�,�%xMIM�.�P��׎#�*����1�"�: |�f\ݿD}��U�lG1T�X�/\]��#;�v0G�u�`��lQ�����=�P��暒U}�7`���3��k�~)>�����J4�[;;d��*����x��ȗ�pvj?� ��+��>����f"�F���Ձ7O������,(F���U�X$�1�[k�C��uRB�J��HњlvN�	k	jp�I��َ��%n�E�W����X��k�D|�B�05�f�1�XL�7��ocҁ�CW`��)�v"dE���};	q��
U�
���R=T��ZVV���V�NE�����0���{���V �����D]��1���+{�9D�U�oޜ�Ɲaii���D�e�k��ˆA��@�i��W��E���������d��1�"��*�>�t>~v��#nm��Ų��r��w�ͥvW��yT����[�X�d�d��bm��IUֹ�����C駱Ԧ�{���FQ�����r����_r'���z�\�tP8m9�زk����^������I�|��)���Ʀ��f�RD�<Y�0�#On��a��e��s�Ͷ���2+�0���B�p��~1��.x��렅���� (<<B
Y�Lv��d��x��$�����Ϟ��S������,��I��T~�䙫e[��u�w�`���Koi^�n�=�����V&�%{t�9�Fƙx�pO�;K�z��[�2�N(w¸�g~s?RA׺:F8�ߔf4S��C�������6��+��k.�L%)y�5��n�拊�����]21M����m���|�  ��g?��{c�a<�# �޻�b�4zzz����N����y�^�����a�kOW��Sd��]�?����|;P[S6��CK�s(�2�Xr,��R��E�^:<�Z�k�5�?�:G9CC�Ap�h�$�^P�q����|g!3x�en ���ݷNvf=	nۊ�,��@=d��v��$������v�%!C�\�B��W�%�r �?�ʃ����<cC`�ƣy\&��v׉e�
B��1�.�#��0'� ��5��#	���x���_�J>���u������#Aq~�,#ŝ�S���g��f&�aJQD~�����#��c���L9��%�<�a�P�Y�s�yyy�����Ż�}U�y���%uM�.�I���w�?ã'k�_�^b��?n��`@oX�8��_�ty�������忮!/U�Uu����n�]l�%$Z�ni�wW�~����+���8�E$d�����I�$=c���3X^�l����a�!$���zF��Ӎ��0��cVIr���#$d�zY5���������$h�=���q������5��;��c� �İ�2V�9�:I۴֝%M-\�0���s&�&����P.��}����Ds������������BA��PP((

��BA��PP((����myh3q�an]�xE=���ҳ"��ErQB�E�X.�k$,��,��-�y�-�za�����6�`⻹oSE�=��ڦm�3��K3�g�y<�ʛM��+W�~���]9;]��PK   �n'Y�7}b  ]  /   images/7f5f08f4-fdda-425c-ad26-fd4aedde5760.png]��PNG

   IHDR   d   3   ai�   	pHYs  N�  N��"��   tEXtSoftware www.inkscape.org��<  �IDATx��\	��Wq����c�{gfgv��5۬/��)F���("�X�+R!"F�����#Aز�m6���]�w�;;;�s��3����w�����O���.�ݖ�7�]��zU��ޫ�^�]���>D��)wb�d�����p8J�M��x�Q��iH�xڇe�3̣��zI��V��ϝX&��\���U�9��:f��h�P���$X�pbf�!oV�+��
h������i&�j�fJ���Q��0��� �97:�bН%)���#F�w����<�%*�V'��z��fs��Qxg:f	��P
5�����i�Iöi���S�o0y�����)�C�����Q��7�{� 3���p��ӄQ�PG�!�U��;�a:�L��	̡�߻�s2�k�2�	�;�����8�eH�<J�Q�"ux�n�`DC&'��`�0\�`�5ޥ@z�, a_V�i�B�=����e����qd|l������E�{:ZW� ��E��{(Ң{��v!f�?Y�������)wsǌ#��q<?�B�%�*����М��B����ᖫV���qz�O�T���L	���&X��^ӖAS��'φ��u5���˵�^�:nqî$��������ݽ	��fI1�M}o��!�v�8�v ����XN�7���1�<�䲻����%0���ଯ���z�486v�3C3��SC!5��jΡ�)�Gτ�1)o���
�}��Q���Od�b�Nʏo`�)�ߦ�eXm�ؘ�.��ߝ$'��F�%�􌏤t=�����6�`��[	�$t"f@��D�If�ҷ���Й��I������^"WXc,!X%�6M#��(��"b�;+�$ac~�c[rK�J���.��?�u�|h38�X��k�R�f���1ˮ�W�c��^Ni&�X.�*نd�K�,AzYU�λK�D�E�
�'=�$uWI/�F�%�ؕ�`)��� ;Bm���:�t������7#}s���D���Ӥ�]�0���ۚ9ƶ��y��ʙbO�g1a��!�b��o�E��I.K+(�ؠ�P�pV"m�M�M�QOjP��2+o��l�4%@ӯ@_�`3�-�dn�k߇���Ͱj���c��H��drVJr4& �t���	�'�u;������Qlܽd���\T�E��P�D#�9�&"��^�	�6U=a��(ڝ��r�Rdx��!���(�</F4j�%�l�g���G��w��[xn��"�V�n�S���,X��1��V�4p���t�&Bv��P�,a��*	n3� �A�4�{�}���y�m�h�#�����(��wt�&Lj,����,����&��6"�/���4�B�p�:[���#3����Cس�C�?ta
��*Zښ���$��S���mGMM~�h`t|K�q�j/�~�&摜]$�;��gjk��,�p��d����#u����1��Z�;��X+}��� �UD��W��u#��`�ܸ_}C#:;��Leqfp��\�����	~�|���R�>�g%���㖲<�2C4|�8�
�Ģ�R%���l��M�%�]�o��d��	��H��Ko�V�5d`]N���ʩ���P���ġ���IֺX,PZ��2Lw�|����@*�&"9*�P���JR����&L����U�A��ԖN�x�j��`�}�v)U��_P�.]G.WRmҏ9T'���ߔ>G��K�_�Z��TFn�p�o�M��ot|Κ� �t*'F������
�h�Q��ф՚��XM��K�Ee�w��9�7=�$�`0�g���<�BmiV��Ό
���C��C�E ��@3��Bx�0>9O�Ε��Y���qJgrg!�2����2S�o�����ĩ��*��R�X���s?���VI�%$��a���vQ�]�Q�l��W~���tn�qc�[����L$�B���-x�bi���� �����N��l ;щELN/m��%1dc*)���'M-��1��b��084����;�N�q��I�����M��>���<�+�&Hsش��%uLل-�V+GL������XZZ�]w���_����'�p:���[m����xu���ɞ�������Z%�����u��O�63���"�m��������ӆ3���'n;�mm�HҶ�c��<r����|5�UV�|m�k�:9!�M/�gf�h�D[��ر��BKf���dd��%���<v6���r��Ѿ��ؠ�B~L�,���w|�3x��1ڳu��u�p���ٶ��,f
;����Rf��[*����,�y��7�=�N݃sS<��������*�F��jIL_�������S�s�\d���=�C��`�LY��>İ�&sCG�_�닸��G������|wC|��{��lY#������S��u̷��3��1C�]�Cf���&Ƹ���?��]�+9��7<C*��$�.�F2M�By��e��/��LF}��9����s�o?�.4ԇ�9��lr�Y?�啛��ێ��%�%Mՙ._U�,�6�ȯg��c�V|ʕSY�T�������(�JkOkR�07V��夻��V�; Q|�t۠�������(��ne�uy�:K~$�����o�:i	g1�⛿�AW�Mi<p��*a��.F�.�ZBg
z��x�/#\X������W/�POL���tgwCڒ���̹_uy�J3�
.�dc����ئU
۔]�)a'.[�����zJ�y��Sg�w�eqxw�4�//���L�d�t�^S�&u���C�꼁w����l�S�P�:����V���|܃唛�*�Huu��S_bWJ�oL��*��ģ���>�V�8�>O�������n��c��ӆ��9!�}��/h��c�rN��li�E׎f?y�޴�ӋXX\�C,���	��I������D"]�������*��thW� a5ľ�;n^�(#��K87�ώ��:� �O3����������o��_�^o�� �M ��������|��9O�L��_�w|���G߇��>bPZ��q�¤����j2#g���`����� O<����0�����<�����u�a2�����MfO�[ɠ��Z���S�g�3r�~����ŗ.���dp䅳��Ղw�z-j�|ph�iF}�� IG{[�̚���i�v2Y�ֆ09� G��\ՅPЏ=�;��{�M7�G��f^A�sYe�g�o�$����h�S7Y����5!>�|�]b+�6̱Cp�������VM��A�0��3���~�� >����} m��8sn���b��S������8���)L.�֫,���R*�Q��b�:1Ad)N�B�ňo؇G�|ѕU\����)Qao��]�z4�u�"���BLȡ���lC1켨���%��.3g��<Bjk�;���݊���T�V]���ZA�/���Gv�3��n��:ë�'|�$:k�djR�=�����f_�x��uV�RM��5�J;l+N�ˌ��3��y�lۈ���Ɍ`f2sy�����I�5��f����u�)�3���o�&vܵw6�=�p�/z�qg��n�^�sn;��XKj���;*�)֗S�e������Z��՗�Nx�{t�5����U�I�����:�d�{�� �E1�LM��e	6_�s_�.���W�L�h���λ������M*]'՜�����ǃ��O�^��
3!�+��<Fj�g�f�`��p�>��>���y��� ���7ϋ�2���5��͠���o	�xjU�d�����u��� �mwh��O�����+���]�;���j�q�����a"�W�Q�R��g���|a�[l�����L}n!Vv�t���k�z$���i�V$2.��mf��VY��Xd�*_T�\m^�jȞ@�&�~&�����m��28;p�--�����S����h)�yѠ���r�U��y+Icf��qo����=Q�U!�Wބ�ZKl�x���ބ��(b�8��owbp` �@ ���Sr�w���jo%��K5��J���ϊ��nI�
�3rE�kz�c]^��$/��Ey/��y11>�CC��|H�i	~��W���Č�]��юK��_cؐwv��ҒB�z%��.�PЇ��y���������;�W�]C����7�n��KM���'�����;W�0艧^Bm����rs��sϡ��7�r���En.^n��b�K�tPn���U�Ea���M��~�-�ު��iټ����M^�b	�������x\�`Ng+��pb�1�NDԫ�-�e<؁�#���'`��m�\N
��3rH�ʤv�k��H����񤱶��v��&5`Xul�z��Y�`��꟫���G�	&/������tխSG�o����m���6e����>�ۉ��4���G�mү�򂊗Y�)�B��+'Fpwo���W�i<w������߅��Z���3Y�85,������\�wp�.q�O�,b|rA}�v�s��%��oO'��=�L���:����?o��}t�h��؜<.�r�!�n/�i��>,���xF^4��r�Į��]��������s�s��ӄ���j���*F��RG��/Z	���=ޗF�u�^d�"��3gǅ��a|��ߧ�[��b�)�Q���(���y���~^eXXYB��Iĭ�|�`���I:�f��+�����D���-={�/,��cZ2�$lq9A,R{%�J*O3o��f��Nb�I��/�^���ȬH3�V�g
>�OpD���.��0F�%-m��T���r<��Ub�z�-�+���g��$p,�[̀{M�E�2�8'��-l3d�	����)�!7R�]�ɁD|	�ļ ����`bb���sI�K�4�#q!�a�h��[o��))ǁ���U���e5妁�H�F(�L@sx�r["6�Ċ������C,�����KF>���*�y���ޟk�o���22Ɉ�a�R��,]�*r!YD<�}����1��>L�1h,��g��D�dB�1ᮤ� �?GDP�+E��H����Vy���R���6n�yЛE{m\�ۨ�.ڿ$J	��9�連)��@$F] %Ag�eeM"�p���`w��8� �)�j���ql���0v�.��l܏�d������.�f��9ڄ��hJ`;ڄو��&8��S4T���`Rpb��,�֗�ߓ�%I``cZ+�E*M�m��J1ֳ�2�8��͕��fH�̢�;�Z�#����q�1b�	qdP�:�!W�Ys�S��80�S6��r�KĔ�Vua.+$�n�@H����J�S�7�'PD�`�DtuH��ƣ>�R�C��� �0��5��T.�х�!�R�M���c1�<u�nn=�Q(2���fB��pq8𘄧AL��Q|�.��7$<��R��M��� a��z�����k�۩�����o�|����l�WgZ�眛�єV����2¤�-�7KOc�.Y�rT9&�N��s�F�2��2��)<p�N��%?�1$��'�T�	�Wc&�N⡗k�-ZoΉ�o#�/�D@�0�����^��-3��p�R�f8�U�9�{_{�F��)���а�9+���p���b`+���ٰ�&�1��ud��S�"�<�0G,�MJt"���@~��^b����jl��J%C>C�����,TȠN�����D��χ�s(��[+�i�d�T���OPqY0V;cKLF��rr�鱁�2�$��	_y���-��,��c*���\PS����G��̡��0�ϯ΅����Ϗ��ݹ�h@چ�G<��S6��YqK@a�5�(1��ӢT��d���OBE`�G���Ǳ!�ɏ,6r���]f��$�ӎ���3D7s�2���G\k%�(G\sav���}������k�f�6����0�;Ov))1�x@���۰:�J���a�r�yC!϶��b�hk �dG���Nd֢ޑ�X*���^�.kE�c��ޱ�d|�g�D�c)ZQ�8��4{,�������L�����a#8�}�t�?��q�d�    IEND�B`�PK   �n'Y腸��� v� /   images/a03bdc4a-b433-4a71-810a-a5f1c0469152.png�eSLЮ	N����ݝE�ww�����tqX�]�.��=�_�z��k�SS��s�P�FA�G���B���P�����?�����6mg((ԡ��/)��PP�������=��&��D�W��(��1�RE"H6"P��(D3�OX(�ſS����~>�|����&�3@��/1GƋJ�/�O�ev�'��Ӻ��j����R��"��B ��?'M��7�GSY��ޗ�M3B|�2�we�� ��?E�����o�-=��.��`�v�I?�P槢��=䯳�?0۬�$g2|�.�T�4+�*0;5C�!����e����|�$SPP���K�C`�:! ��e��q�U:������4S���Ҟ@�߫���Z4^K�r�t�=�ܖ�j�~|E�"��D��X��2��h��-4S�lW�W�����6��̊(și�����,�.X��Mų��ܑ�EfEک��C�����^-�ܺ=GOeyYZ��VS!U��>dc�b{�h���ԕ����/��<�*=+bef�����VD-��޷½wj+N��?�����aK��4�鳣�OLtY��H��O���'\�������?���y���Ny���~g��TZ����W�w��%
=��$G�M�����Yl�*�e�kgwL�\����)���p>�����y���4��W���Z8b8@S�磏�S%F��V�BsE��bC�zئ�:�T-�j�R*�8���oo2~���}lt���d�[�u�nYo�q?���ܝ	5�����.��� #s4�/�d���RY����V�z_2�G�Z>������d�!�fX�֦��ئ�sɱԮ(r,.�abj��({
c)sP����f�:%U~ɸ9:�B��s(�o�����rvZfĔ���vX��VkT��h���f�	�؃~�`�����������-�t�qg]]5���G
}\䟪w�0$x�Ф��-����Swy{>��,丶[���l�.Y�V �up�'�w���{�E�	�b��[�LfFaB�U�]���Julގ��]�75�Z3��U����?��z�E�-mLa�����dN���Mg�3W4��y�����*�Y�e�r����:�,�A�*��c�4L�kr�_~�4�ɬ��~Kc�/˞��r!���E\�O.3���q���C�M��H;~I-ը�$%�����Cz>E�bf�K�$0���+�t�]wA�*ٰuQ!��*�����3����8�ș4׆�e<3~��ی���;J�ϟ4j4�����>���[��%���:7�[{/�����(9G ��Sd�n{�sSA��1����~j=��9�1��C~yG<�RTr.�)P�.7O�)�U�)u���8[�1�2��_�P�d�
=r��n�F&8a� �"�@ :s�AF���dj��
��V�G�����p��� 1?0W�@�oX�d��]��s�KЎ������zQ��$z�w�;����P��#��X3}T���;N��;�8x�6fu5�~F*��Z��e�x�>�!��o� +2�˩�0Fô|#G�/�J3�����Y���o(��j��I9�N�d�7��k/�X�M�����8��[��J���_��uuuS~����J�,Аy���������:.�D�7f/f�dh�M--/ۭ�]<<G�]���e��n_<yu�4�i�o�&_{7����s)�q�"+�U�ݐ|�z���1�E��Bē��y�'���0�/}:,D�;�b��ع���呂W�=�O���#ːn�R
4@u�<��V�$�6�)����K7t���(��7Wx����:c���?���j�R&�r����c�r���B�%W��|O`��ɰ�����0�ǓI��_�����c�N���mc� �R!�9����9�⮃��l0)��z%���A�Mq�9_��h��TI��J�&%��0J�����Q�f��A�+hV/�Z�@M����Ԝ�uR3@P��6[������G�4�$�[�P<�0Ã\avjbE�Ҍ�����^;
:gR���.�@���,��qRR��:T蟙i8[qa!�g����Anad݋�����S>��Fx4��;��E?�5��=����}'�"O�E�:��]��َ+�K
�qZz~LMK�K�};T���r�y�����y}�$��w���f񅇨�2���5�\M�'�薳��mF�Tb�d�#�Qq>�Î;�(�j�G���U��k��?+�\;��P�q��t�$R�5�W����N���L�&�.qVl�p۹���M�7�ҋf�	��A���+Hy5灚�Y���,ݗ\l�G+�eN��]��N�,���N[�X�(�u,�[�@�?���f����I����d�]'2kKy��Z�FX��r�x�U: 1�h���,� �2@,-@7�0I�9�K_�q�>�ϝj}�?Y�Y���!#Y�\v<����3��%O=Pf?��e��PL��Y��5�EP�m�F9�1��V����sR�P?Q�G�3��!: %O�3�2K�q�;���R�I�H�>��ߦ_=,�<L/}x��.3�,�=�l�V.U-*�,�q�ĳ�6Nج���L,��pu��q_w
�:�� ���E	�,80��"����G��z���P��ՃIA�`�<U��s�f;P��eX��
tl��N]�Ք�j�~����b�\-�,YQ�|?:� �0^0=5�1�b����`����u�e���!f�i���^4s*�t�UgJ�0F��g�gy�O���p�=��+>��R�_�Hՙ{- U��������6����w3�+1Q~4fI��
-0C�����h���A�a�B� m!g��`M-��\B>r`�F�s��g|\���L�a���{�[Q��ѩ[��j�}�`�^����0��SAb�.�P2E)�Tz�<��8���"Sd7P���hdx2�����dd�3Y��`H)�D�����I�<�J5l��*M}��\K�9�@l����s#�>�V��D4.ZUh��P�/v� MK�B��4F��Sl�����������d�_��v�Gx��6����W�pm�y�b��8�|�͟':䎞6���^i�C!0r��#���͆ؒ{�_���\�,G�s��&�o��^c��<UÁF-�d���e%�T���t�W����(���Q���͏o�z��9���N�ܵdqC׀�'5n�z�>ν�_��|B��� I��3ʲbb{�"�P���6Z[>WKk����f�}��co��/r�ɫꢁ�ѕ�)x�	�Lg��
�9(��O��J@�
*��%):V��
G`��i��_�1���@#U��rmMJk )�V�b�F �<ލ<|�h�xZ�q<�!HE�J��K)����T�{"��1�jUm�_u��q��`e"a��#i[��P7o�͠�fB"f��CU����x����n�W�]-�V�U�4��nKF6���)e,���s�H("�Q=������y��lQrC�ìP��x����/v� �p����B��ߏq����
�.�}dj5��LĬ�	�2�"��z���Iݓ��[����96�1J#��#�Q+����YÕd˔�[8���"�h�\���l�V��X_�
��oҶ��ҕ̺�� �a�W=�KYu}{�~����Թw�a���������x�1(2�[�3W�۝�'�@Uq��J����W	V�#�_�>��0�ل��0��·���
,�_0Y�h �~DL8�S`5D5bx-5UDq�]g���=�l�Fp�� ��F�u|�6f�iU6��z�"��7C���4:fx�4t
h��Ι��y�Q�',b.xn�Z�4ш ]0�h�^�|��1A�'\�5CR��6;��sS�:
�Fd�Ј�A�R(����}<�?�������G.F*K�n�o��o���<�t�%cw,DWH�Y� �J�UZ��r�����Ԯ��-��ަ3=�ÎE�̀��L�CY2�`�{>�D�Vr��x>�[�i�Y��_��YY�� \�BX�/)ڋ��榭">B\$T�).����"���:W��@��>��t.�4,V����\�.ךw�;�k͉�{��{�q�}xe`�2����G���z0��m���"��}� m��~�|%¤����+r�~�^ﶾ�5��s��������W�$p�#�B�_[�x��d"2};�I���w
� -�l�o� ��l����Zl�,ϓ��t��r��= K�b0�ȃ����{2�l4��7�j�LLҩ\�2j �\?#l=�5����C">�����f
kLH�xt���Q���4l�P̀^C'���5L��|��`��e�r��`�H�۔�MB��-ǔL#��,J~�t�Ձ�j�N�O���[�Q�~����z�9�'f���L]��
� ����""�:Y%��qd���.TM�u9G1�oi�]{2_��	Ew=�����Ig�TD�ҙ �X6(��������MV��OҚ�Z$�/�<並۷x�N?z��2���9����k��a�=Κ6[Á��J�?0�5�?i_����g���KO9;�ͪ����p|��soy<���}\p�=Oirqs����"G��n�Kx����*�y�h6�_\�q�0�]�\"龹G�v�w�tz�e�g��S���'-�I�i05\H���͒~9Y"� .��E�0}��(��G�A��"4��UH�4�?�̗�����r�$F��ƿ`��%��+������ƒU�~�gyT�Y�k�+�I�WF���bXU��ґ�Ԍ��239#܏�-b����h`��C+��́��bS7<�TM�I��~�j�V-��8{��P[:�ŐB������h�R��� ��6�q@�����W@F�NNf5����I�z���J��(L7�h�5�V��2��-�P��x�k4�0�X���q���|a��C-����|y�H��#֬!��5��{g��Xw�-R��cFC��5括�a�m.���}헊�Z8ovL\��ꤾ<伒fgg���n�I�]@t��=v�������z{'ɧ\�i�^�@���V~�H����c���U���6l�f�wy�������i��x���*#����ު�\����z�d/u�=u�#�4{�l���%"�RRV�&��G�j��Z�ǯ.��W�Y0�N|��*���	�
M&�¯�y��R��,2ER��=�tQ�9��ꈚ��E`x���r	~gju�!�u�n|mW� ���a��v2�����ү��Zm�)7g�5���eA{3˵ǋ UuOB���r�L��Lj%��-=���Sم�E��,v�!��S���>X����C�,�X\t�ֺ��}dJf����t�$�������8���Qt&�vv�����\�^�z1�_n��7��10y��75*g�?ռ�Q��m�R5[�x�!0�m�p�. @�cr����!���!p�RO�a�2�$X���"�9�K���h}�8��h6�xRXi-��VLˎ@�����SDA;�0u;�����|Sÿ`ɹu�v����Ƭ�7.�І����;�]ɕk˃?*/[�.�j�����m���I��sW�?�#m�E��1����۳L�"5ex������&L��`�����f�/9B�;�V�?!�ٰ�%�>�u'D�$ ��#w��-5���C�a�AT}1�nsM�r�����C�h'\4�ņ3���k�)/�<.���?�P������9�9,���N^���	�nrf��irX"J�B�2��ȹ��v�E����$��,��,'���� ��΋�����e��qg����s��4J���w�g��������F���� or��Ns���qz��Jvog���2�����J��5|ag����`���[9������mT�-΃u&��z�V��5Z.k�n�4�Q�Ξ=3:��o�7�.�f�R���V�"lV��!��Ђa-�Yv W�HCa�M��%�}���$2���N�ќ+<��9k�	oں������E���PDt>7���`�H��y�w��gJkd�̰�َlk"y1����f�XdlA�ț�s��Rm��F�9�F��@Q� b����^[eɚ�ޜ��4q_���7y�xۃTJ˼�p�$N��r����.:���W��O������L��5.���nG�	��n��n޻}ܭ��ú}��IQ�ة�W�u���K?�[*v\�o%�}�
�����(2��<��WY������t
×����������'lJDb���)�dτ���h��j>z�������=�9���P���_�e��.hr���˲�HN�rh����r�H�G%N7*���Ŗ�^-�����m�y���o���IM��y���xl8��m���wui,7R�o*�-�#�Oc
��¼x2�����l��M���M�J<S�E�f,N�L����} ����b�Y��8��-�B3�����x�߳{lX|�(�Q�
�c�K��8�s�-7u�ʊ��o�L��9�K0��Io�JѦ�g�Nl�i��x�L歐.r��kY�.��;N�+�8��4�'j�
3�BX�{��W��0F$5��(6�F)%'�,H�1٬G����m�%��<g�v��u������Zk,��h��u䨃T�խK3P����kzK�$o����zޫ4��J_����ݼ��rṄ��2<�hTY��4��o������nv*�}����
p{��:;�X��C\�dn��ޗ֩b�>�C�_�.k�)(�(�"�t6�G�;�<ŕ�9�8$�Z����9�6� ,g}������T!�� �'
w����t�~�	UZCC��Ł��s�
�����㥯�����>�0S�KY{w�+12c�Ҹ(K�ab*��z���KxV�JQ����1<Wl	��6iv��oFe
Q��<L}�N��42<z3�S`����_�m�c��4������Ņ&��tϭ�g�<���a7���V�(�T�h���d.)����^X��B�lj�o����ũ�:�;G_�4�W_f�5u��d��J^� *�#n;��i��4ZC��p�A*r��y�x�k�NX��|XY9�feL9}��=�)�)�4f���+�w�h�*ځ�I���h+��q����k�Z�����P�-��]��F��ˀ��ڪ���c�7ܦ�:=W8K���~��l�����Y7�;5u:�������3���\����IO��t&P3k	��	Ȅ��t���JK��I�G�yOC�Q�J4J�Clg������j�=�z����M�kY���!ǎ�nH}=��S��؝��<�zz�M-�#NA�d�j�Vp�����vY�h��b�2�;\�\��T"�\7���m�=����h��Sݑ�7E����*G
����¼����bgG$��.�!��j��Gbl�O�^==+�U�Oѭ�a��Y�����BG�u��Єzj�}�*(O�
�d�6D�n��|�� Ç'�J�4�%�x=�N����M��-Zb�T[6�_4/b}U@�G*�ů�~�u�����'^�i�,��̓��"��`F?�7I�lk�#��̩���G��Ƣd����.���|��B�2�9ck�V&�$�d�l��rryi�nNͧ��|/eɰ���:����e/��� ����w'�CS~iz^�6����\%Дj �<��u�����'���������[�j}�ғ�:E������\Y z���ݘy(�5��n[��)��w�c��v���I\�*���*��.fd��{�&z�[�R����fJO'	��D���?sү�������oO(A]y�����5��[�+>mAu�5K?�^�K��4����<��1���oL(;�iIM�M7���������O�T����]�%����:�?��<�?����tP�N�y�%]����q��I+���xI1|�x��~!ҙ<2��\������g��e�v��i��{sT�$!Pv&�e�<�x�/y4�YĘ����ZF�h�p���ᒷ�Ͱ]�.n�qu�p�K�/�JS��c�����w{r2�7��@ʤ�� �ڜ��k?5
4���H�]��:i�m6'76�q�3:�5s%��C��j��Z*M0%VN9P,i��E���V7B2
�e1:�O�G�\3�<��,���Y�-F-i����U�o�Rmv�����sW��	  6�ՒD�	_ɺ�x�^T)��=7Z5\]m��$h.�CG�QO��W��uXO6���g.C�C���{>]���Rz�J���ZM�����׍�����9)�/�Ey���!��� G�IAj~�G{6���/mf��ۆ/5�Y��Ejo��v��jl�h+�h�KQ��м�X��M���C4q_��
+�g!+�ŷ��'Ζ �:e˵B�myĨ5S�k��|�Ι>�;�_�[�n�~�nx����� �������Ӕ��W����[0�4�2
_��Wϙ&-�[�Z"=,R�m,�5ǧ,e��-��J��\c�w�7����c��EA���w�'ymlM�]վ�F��{��.�ݱ铆45_�[�+�����b^Ԫ��T��2c��d�-��=Z���ϴ�s.����aR9G$���r�������ِ[o���6��Dٻ��b�x����J�e���������!�;��{i�h��?��m��2m�;�KGp{��>���T�Si��+���;��-�>��!(�4d�=M����VTL��{���wW��(DUӌK-��X�1Gi[N�2Ԓ9.=|��Y�~ozi%-�:^�	�B�Y�mmi�Bp��Tzq��B��<k�5���@�fx�U3�*21m�E�@���@����t�z��J��L{�@RU/\A�"<�1F��`t�k~����|x^�> ��2�3E�'��S#��ӵ���F�����?��余8�V����(;z~��X�0�G��Y��b�k�l�EPZ>�E�XC'6�"b5��Df��=6������ GNE5')�A��86UP��:�- �^�a;�̠*����P=�����Vt(�
�-�9��fE`ݚ�V�H��]�r��\=��}g?�������Y�1~�Ѩ����@&�d�����|r��Z�W3�@��$2BrC���QÓ�'_�#��[���%P�����YaD��I��u�[�����T0/�=�E˯V׊�r36"�����Y�%�J�#��T|Y�>/��r��O�L�G���*&����S�ϓ݉�~�e�����1l�[�ی������D\���?Bd�~ �i�K[�+n+c���69a������8��{�|^4>5U�C}8�n2��^J-5A�I�1�c��?f��O��~�=�wq�8��[b�M���x*!]EMf��E�C�|��>O��/pZ,"���ڤm���PF��fk��B��ݼ�g//a�X��P���OQ<-xj��[�
9鱍�D����0���?w�5����vD��Y�:��!��[����Xe�vӿ��fV5�! τ�����8O���s׮�ɨ��H#=a���d@�r�+��$	���}h�{�I>��*`�tt���zx9��3�྽��^#�r���G�K�E�V��Ɲ@pRU��A.E%:���dP_w�q�jD�����%���I�6U#kJ���7%�.5A4mF�rr�h��K�� .La"�Jq*� ��:��KoQA"�PвQ���ĄZ�S � ��.UU�Z����uJ� 0z��������޻86|�q��ش:GN��~ʹwu����|�K�*�r�Aj��K˵^����lݴ|�[7Ĥ&����%8� Q�H����h��|ڝ�6�[(�{0������`�D�u�e��:Hv�\i� ��ۨ�'*�I�O\:@��P��{R:��Oy �Ѷ�CSVAa����fպ�=H.��w�MNp����_w��~��_:Zǿz��ڤ�è����C�0˪~�1�C�x���HJ�#��l��}.�O��y�W�����w���
;��\3���Ρn�@W�I3���2��u�'PE�=�:Մܘ�Y���{��6�U��>B������z>�Ѩ�K�i�>�zb�{o�5�x�H� 8n�?&�+`�#�{87�k;�%2�c*-�^��C<	�"���`w�~m�B���LU=�^�f��;�bS�p��Ԗ0(��-���Dm}�>�����A$�+�i�͓A���ٍ����:�_Q%�&�'�{?n_�8 ������{2�� �]D�F�~1@�y=�]1��X);����Y� �����aj������G�A3��u�w���J;�d]�'�9�¥���@)���c��S���e�V�L���]����3s�3#����*�N�Vn9�fK��ŗ�i7!�,�֙�qB�6�M�x\�da!�R%�kE�-�*Bud3��r���â�}�?��O�:���j��d�U���"sL+_H��ɉ��L�0�_���WmG
�T`��?��SB� a3mt^A�� ���Kd�>s4>��̪Y/�;�g��O0�����f�\U2F*�x��+�N���6�\ž}��<�$�(��$Ghr~{)�m��g���@!x���Y3f���JE����ڶn�S���Qh��Gu	����~�58z�\��x�r���y��?Rj4�C�_[YY(��-��|cZƛG�B���b�b����ϳ��}'��N$�
J�An�e}%ؕ��u ;�)���֥��x�V�*ڣ�+��?#6���)�X�#�:���6d�q��z��-�4 �[�3�7�$�di#�*�����c�(R��؁[��H$fRD�9	t���Sv�2m&DS��Q��Ξ�(���H��@����-a^��#I���`���P�]	���9CS�}6�EKU�؊��!���G ��V�۞����������B�S>.f�O8�]{71L��z}x�s{�tAY�7��(��Z/��2���y>Fw�2ʆ��y����%��o�Q�kk|��<�]�&��?�M�=�(-s�w���*.(�M��bþ��%LG���9���l{�l+FT��҂���2穆�w\��iT�����|�oM�r�xE��^8+����=�uC������o.��>���ʲP�!�����%=�"�s�q���ݿ����̙$  �ԶIf���_�el�8ŨU��mm#u�Wv�� d���OP�7���F�Nv �&���P�
��Z�I��5I���'׌��kQ�����	����Y��i-aJ�w�FT�S،v@�A����'U�I��%7Y~��{k*��L3�ҹ)^zg/��ѩ[Ɓ�e��Fj6�V3j�� �z;�r�~��T���V���D���A^���o�w�9$��e�ŏ{���i-�nâ`�_p��<p�'��1��u�����e�s6��Q�2D��M^�|�EG����6x��N
j�;�gz�y�r�RTP�;Tg��|zͩ�ɹ�=��-�����Wk��Lg�R��3 ��PW3�d����cb�ª ��Q�S[��z���lyvpml~��}6��=�D~�㗡 �hZ���<��&@�oP��w�Վ��WU�P}S���>b�i���tT%V��3�(9�nmS��ʙ��#Z���sN�G�͝MW2/s��y��m&�(� I��S`��ehNm��z֞3�A+�1�n���i��Aa�Dr�QF��_�[AVN	0"�n�"�izᐖӏ�!O �G�^�z�ڬ��3�6-��~�����8��~�T�:���WR��[���}[�΀)�_g�����z��G�z��	M(��I?s�Sh����j�8����q
��`�n��v��렰�2�BE!$t�q�kJ��2�}.�a���V�������f��ʿ�z0�x�w�����ܓt����`���E7�Ĝ��w���˱��J{��Lt��A!'Y�����c��K1s��S�M��Q�@�zbov(H*�+�,�Ggڦx����7M {��/��%�[��ߝ\Rݿ���F��8�\
��)�,���W�����\��e�4�r�(D��R����f��VI�V��r �����
7��˫�^��yAL��V|M�r0#�֖�[_w��/�"�Jc��S���G����N<֢�~��y9�^����`����@��IY�1��/�`�fɑh�ǽ��[%v����ފ�v�O�俴+Ҏ>��ԋ�Rbk�|���4f��h����)ĉĠ�Vb8_��#.Zѝ���'
'��hE�í���� z�G�S9z埦#�E�@�ZAā� ����#L��w�)Y�����IΚ������3ԕ:����WU���V�=�9�I�)�6��k�0�ȱ�C]-��x���6Z�}aM%�^�Jn@Ỗ��	ԥ������/����톰y��A���������|%�ݯ�b�c�:OSl?)P�2Ͷ�Q�5��R�D���Ÿ�	��<�4��>�Wa� E,�mw�~�pi��ɶ�-PP�2H9��:H��v1�ۑ�+9^�L���h���ㄛDO�0�xk�chD9)H*%�p��/�Y����ל��j>�uD�Y����:���@�	���8�D5�,�JÙ�B�#�;�N����9t_I��v�����/��4�t���7��Gz�@�I���*�UӀ��9� )P��6�_=3g~uG;l�i$��������õg8^8��n�IᨓB8o`�*�z>�R��Y���{q���N��r�t��EDb_��f�HВ�4gî`�;�x���s�-X~�U�}��Q��>'~�� �C�S��ü�!#�=Ű�ó��P��c����}U����L��B�5~H-$�6:��b+n�,!�������,�HMM�9���������I�!���&V�_� ��+�2W��j��� NW~T5(�o�0��؛��|��5p���L2���Ѫ]Ϊ���\�7DA�]�͜�p�����=��ܼ�۝h���ݞI#�'H�=/tD/�!���E�NG%���P3���y�⮡����c/k�	�i$�:F��Ղ;�~6S��+�QfB9ex�����ʷ��wiZ�P����+�H�l���6TPa]B�%���ބ'򜛮�{�`OH\�[���1��p%�D?R�O���q�}b�<�OC;�t�P8�q������p�]㸆�f��M�Q�WN^Q|��_�t�q����ٓ����^h��T�N���ܛm�O���n:c�n�[������n���G��7�<��ߕ��9�}��[[ț�[���[a�$8�O8��Us��j�Q�
��y	���+äOы^��^�Eв�4b�`�-�ӄJ�	A�?R�=n�f�zΥ�d{��nN�m�0כPR��'O�㱥�4{?��N{���[n�V�i	���B���Wϓ5 A�.H$,L@�?��X���چ�+ ���ۑ�cl��R�gg&��p�d2��>�~DA��s�~Keu6у��$�v3e�~Ҷ\>j�O�gof� �*�Q�bV	�_S���s��`H�L���L�E��Yk��Τ94C~`�z�6�Pͱ��QdO %X�{�#'�ݜS.2<d�:���Z�9���	V7�Xֆ8�s<�8�kC���4��3J�)U�4�~� ���ѓL~C�R��И9Hն�L9v-u/[-�n�1�.��j��1k*��0�d��"="��Aޞ./���a�P`�Q+zz��j$��#B���5��?��\�/�J�'�I|�����	.>:��G\�92�ا6��bC��ׄ������wI���"�8P5�Q5G������n��j\V����
�&Ψu�n��+�P1����j���"28�(v��~;NX���V�C��zඞ�ۅ���:���8V�M�-�U�y:+p}z���u0 ��sI��/T<N�_)��xּz�X��R�V>����?����)���jE����WT�TvJ-���� ��]\��֠�%���~������Z#�mߴ���;��ʆ�� �fP$�?	�� ��-�ѧ�.�l�)Q A�]ͣ�z�]�>���X�+����Wmb�f" �5��@ݩ� F�"1>��U����c\6�tJX�Y�39�w�RF�Y�?�Gq�89������c0���[u:=�nm!�p���X��o���߬�8˔8�+��J.@q�^��ʋ��s���><��8��$���Λ3�3DH �3z��!JA��)q��GT�-��EĒy񰲽0۸`��_���!�XL+!���ۢ�W�߅G�޹��ӟD����}��u���:{j�u!����]��<��q�'	�L�~�B�=iR�@:臠z�#����U3�8�{SNC2��W[�b$[���� *w�� ���#��{kK�{vf���H�5e�[w�I�q�N��oD9΍D����<�
�&d�}�0�ڂmè:����(0�?��,���m���T�<~�)jC;�}��Q[f�`V�����=�czk����m8���,�xd�Ь� �� �N�0���֬>`���|�
O��h�3�;np��G�?eG=v���m���;�Щ$�9��'	p�
�ˌjtcdy��SX�m�y~ I�}�%�V�x����8�Y'������9J�n]}����3Ko^U��m��eLz�}�a��{Q3��Kg����	����n��bA�R찓��e�8��^<�'Q^,����Yj���s(D�~'-,�&x�E��8�l���G�T��w�-�\�J��0�����K$jI�@}�ŭB��쒙��7�+��ƶz�����. ��h��.�Pk���_@ޢf�p�E!&i�^4��i�<P,;ؐ*�Qa���(�1�8'\?��&�{ }��}�sM_7D�'6k�\B{��î�X�	��C�|���
�:9����A�!�O�!bZ�h�X|���t�	(W/	�����y
����U���@ʶZtRJs4�
��5rD�Wҋ!��}�����Ƌ\��r�D��>�m��Dƒ���X��y�0 �vǄ�I@8j?���t[+������&L���%i� Qo.�
�}��x�0V�K��T��1U^}�3v�ɘ��zX�����	��-^�7d7��J��$Ǭ|*p
��B��caXͦ�s��I�Ҧ���E;K���*<�=���]���'��s�Y���
.��[��Yޘ�ٯ�����/Un�xs]��>�o;`f]��#�.���m�4Ɗ�(m�^�������mx�ǜ�W��>�`�a�;��iǍ��Ϩy�ρ���ޞ���ʲU�Z�F��"�Zl���0F�D�����/���sS�\7��cXS+��5ծx2�\�(?��d\�P.�d�� �\���CD�<4�B�$�H�!��*��7�<���:نYz([�6�,�@AQ'i�ZPȔaC��5-��xSx��=~Z��*{���K���μ"��H�;<TQx��o�JQ#��.���H��U:�T�l6���>�(�9�_���~����n�zd݊~6�86��R��ԸiV��W�@� ݀�&����12'<G��#˟��_�M���eW�1��F���o�T��E!Z�q�u?_��2kB-Y��й�,۾s=��O����'��OYY�H���5U�l��w�}J�_��#WG��)�elk���+fi�2��=W�|�;�ʚ����k<ԾL���98^����!��u��*C]�ـiFZ�`���$�H�&7o^�/=0-�|�(���X�����,o�Q�9V����U�N���5qj���d�I���]�$��:Z����)��S^��r|�\�e�vb&������E��KA�l;[V�I������dk�m�w7c��v����_��7�tɻS�f��7�Z�!��cY�eQ#��i0��(��У�$�v��Q:k4��ҖTY�=��+���6��W�,*}��X�$C�LR������(T��(|M6�M~ԛ�[�H2hc���b���KG��C"C����Ke�a��j����V�����Ԣkn!V��?xߍt�>��>u�]6(ً�P��`�a��e���G��_(0��$ ź`e�:�#��
)�R��D;�'W��q�90��b&8n���:"��Z-jA���h��o���4߯Y�;��N��ս��R�J���3� �����j7�Y0X�/m4c�����{�S���� @����������|Vy~gH����bZO���S���O�X�F����ܾ}��[oS_7z5�9�7��4S��xa�XՕ��r��j��u���xm+�qV�&'��Ӕ�'½"�H�*ד]-FN�Y�UQ!��`��g�)�AMO��$٪B~˱Ai�AflLy�nc2
9j*���4'̚0�PK�+���	�]c�!�F���sq���[]��"�6�*�Mͮ���EXS�.g^Z�5�9ĭ���M�9�LɅ���'6d�,���C��`��:���EQ�)O���i��Z�1�lm�nn�����n�s�:�ol^�w76���3���ʹ�D�W�q�ѿ�C�/>2;>�]�����"<������u�i��l�Ho��KV�-&Kj�v鏾��&���ۄ2���~���'���t|"��}��R���pD�����r@��W�ݽ��VN�4O=bE���%��rވ��DIE�/Vk�V�oU�ȸ�e(�M�k}�h��{�Cѵ���"����8��J�C���� �e �C���)�l%ޞI��<��m�����7 }@��jH��I5�C��ZJ�"���K*T�]�n�t���8֔��5��ssEVV]m�,�*O���P��W �y_ko�ho��m�)�PvJ����h������ۤ��Qp>��)�K!�UN�J-��;����bl��}�V�,�qw�OU$"��W��h�i��,�hW�-;���^q� �Mn_����yI<`@��1p�گ�C��}q�bu����7x�e�@D���s�x<Y�C��/Kܷ<��d��כ��hS��T*0z��`�ͳK(γ�ET�"z�6��-��_�wtP3�pw���������D��eX���)��}��*^Q[eY8Z	Yq�\�N�|�j�[B�_����?��c���H�5�^�cK�9:�yP�'S
���\�ֳ�B���"��
bQ�UV����a�L۱��n�����!H�S>y5�*ٚ����y��H�����ؗ�UbL1BG��T����̪��S�9�콲#�j1~��i.�y���Y����l-�$�PB�%�2�F͡�l5-&�1�8��oxN�aeC�;b��&i8��C���d5��2~���ܨa�J,W��ò��Z"��\٩��,_-���~�*�Fg��N�Z-T���]��u �(����<���X�d����$N\י�y>��v&�߸��ʢ�;�[^�>��/2�Hv�]l���k�6�3D��go���W��e���	�s���}���FI�<�4�~���W�g�KGc�Հ+���+�(� �[w��]|��]�M�m��"M�m�"���i�!����w��ν�Ӱ`A��+{��k�'1ei%�5���+�ER�_w�1ߺ8�f壂��1�M��qL�g�轗/��>�+YV�}�������d���l����Ԭ�"������!���=�PլCY�����9�O���$Y%��x���M�A{�/AN���	/(���H�F�$�	�V�cW�5��{��W�D�D�33Y1AV�=~�_p<xm�0_�ϬvqW�L�[܇��CV����r�?v��DL9�
#<�L8֊��6����S���y�����E6�b(z�%�D��3�^N=Ϣ�;�<o�\��BL����8�B�Je��+v��t:\_�E��9��a�b�<
[��[���E���=�A?�s]K13DD\��Q`Sk�R�\C�f��i�G���[�?�(t��Z���?���oΫ�+����c��	���=��lN�y@���o2������p�;F�w��;������8��px�Rq��1�*[&̕�`	5���;܄禁�4�r>��B�O�V+�h�}�H��d�z��Q�F�1G&K9����`E�6�	�Q&F�m&`�U&����i~��\Ɯ�q�=⹵<����帱�\U����8���<�R�#K{5�Ó�xI(KZM�)VI�͡z\��?>�����9ldKA�� �p
C��*��Q���FB�|�b1����A�v��Q�a��j�~�7޸^�ۙ����n�m9w����������nj8N��hpE�Z�¿	�=6~�K/�NN~6�aퟘ��F��!C��$�h/�ݾHnmG�/N�˂�.]�L7��-�w@��n�E�6��x:JH��+�.��RL���P��,3Ap샊��ZMgIA�$Z�*�>�����j[+R�hK���ΗN;_�Ty5(}u��\0ƚ#1�d��0��~�����*j2�S}c�|\sӍ����@�\p�3z�Y���Td�g�351>��0�/Bծ��]�%��u
�X�Q?L�P[b|�A�e"� �
�)�����"\�w�Wk�{	]^�O+g}��1���I��J�r(;�����*d��Og�����'�-N��C/�֜�p��~�%t�7g��NV�v1C�P�C0�BǸ�L��9����ٓe�q'�g?w_k���46�D��H#ɴ<҄C����zrȡ'���~��/�7�߽�Þ�c{�0GCQE� b���og?����;�nU�A����bu���s�����_��t��p\(��T�De�*�{���9D�����9�l�����-~x�}�|T��"�����<�kU$�j��a�H��a�F� c��Y���:��i������k���\8Z�5U��#���2^�����o;E����og��8�������Ͼ��h�<��|�Ď����_�zL�5�I��Dk�2E���N��Fk2V�,b����޶y;�������e�����qȿ�s�T;�M6� @:88hu:�=�����z�ۗ:�V��쥝C��P+����*�b4������B�R&�Hh�`㊚-?�;��m-8��+�C��݌�}029�4��3�+G�"q~,Ґ3���ٕl�0cհ}�=k9� ��E!lJG�P1��?"�T��%
=��ԃ��)���d�e)e �����RL�	�,�=�����C-V��]����_9��:S>W���ڪ�n;�ƪS:5b��g[[~Q�T&��)��X[������n��s�ﾻ�&���3v#��ECFI�d�&#lH��Wd4 z1<����}��g2� A�p0��;Bb�$|G��*�~/�L�D��Y*XB|��R�5��m��L�-�{/ّ!����bޯB����78vFL9�69h�R����1�����̆g|�=p��{�!Fk�������tڂ�є�q@'��~���O���}B�~_�38�4�7`�K�
Ja�MΎ��iuҾLЫR0��(] ��eI�KG�#UFL�o4CD>�ha�!� ��-B���$�����D��K�s}���k�_�0��Z2�͍63�A$ݛ;��u=8�D}BJ����!N�>�����*��,���u��A�jg�q`�t'`�-�039��Na��L���f�S�7|���Dy��v�,�����Ǵ�ߦ��3	�l>��dL�|�@��	\CJ�깺MI�6��?�)8`
hΨ���[�R����l�|:;���׻�����mㄞ��S��9��9�A�T��J��>�n��RTa���y�w�]H+ib������,r6���8�7�xQ���O�D����|Q�kwh������^W�Δ���Tf
}��L$-jC#vN6ob�l�v���:zV�p$�#I?�S�=޴�#H�!4�!���	�(��@�B��k��nz�6r���5�QF���r͜�z�_�P#�D��L�ɴXE$�9Ps%ӘМ/8D�QlL�E���h�+�n�3T0jx���ش[S�0�=��y��.�����pV��c�ډ��4��?��/a���wr���c0z/�̭���v�hf5�4cc��JVسH����^ΨŠf�Fm��}�C1b�Fzw����H� ��m�I9�-` ˠ\��������k�
�2���c�����Kq[e/���%����=L�1"~�9=�4�W��8R��7�P`��foB�Õ,D'BF�m6�pA	�0~gG�'$>�����pIs2�#�U"�-C959ȃ��{�KE�K����@3U4�V�d���T��1�K6'/63j��Yha��Tͺ02iyT��&��Mv@`�az���>�-K)�I�
��P%*io��I���l��mo4���*�)p�Yy�ŧX�uh�������`�/��p���E�F�v�Ǳ:�S�c9=�َ�S�XIip~�v�vz�}9=;&�]�2/�+;�)hwr�,�AHՓb.i�f.!�V�'�`����w���Η�╭9=��r������7IK_~��-��g����7�N��J��g�{eH����L�s�R����QG�	��|"I�y�� S�6׿��P{wg�·7�nX�Uh�"�5N%��U���D�cn����0���OMqt@�~w�~4R��#ڿAc��ؙ֚mZ��i�{"8� ���R'��c4Ьp��uh%(4��E�M����R����&;�}���j����g
	u�	��E ����
��b<Ĺʗ�4�s���4�#Z���eOL3�Xfv�Ѭ�|߹_�Ն�fs��v�mߏ]��lmy1N�G�TȾu�ܙ?�$5�G�j���Y�q��N�j�9���\�Z�|^W�Y���/�ƳS���^c$wN��#�x{��*4��R�����+���;���< ���4��d�BkX���)A�rFb`�co8Z[M�KP][��_�Kb�B��W��f$�U�-��ڶR���,�,��D
0�}~��\v�Kvakk[��@��阖I]��L��CȄh�d4��HЪ`���ҤracL=���b_t�����[��x4 /����9���vNP�-�t"rc���T �N��h�B@,���B��ہL�	��!0#�y���3���)�t�k��y�/t����j;v5J`|���j���^��uj�+�+���S��h�����Dϕi�4c�~���x2c��d!u��@�\�-��Z�h��&�L�ϕ�f3��,�n{�~�I�%/1��~fXo������U�@�����\�����Ǜ1̳����uZ�Wہ>��{�ƺ��S�.��U���Z�����6
6x��3����}����y����U�w���"Ns�w�Z�j��+rS���BQ�Qτڒ�Q�7-��ܔ(w����a�HZp�F�Ic�o�`�ϖR{M�ߘ�iViT@Ri�ȶS'��h��9rj�|.��a+v�}Q��5[l~��h̟mI:�A�E)��>�"s,+Nc���U*�x6Z��Z��ٯEQ:i��N���Cϲ�{[[pGv���*����N�4���S������ѭ7����|y�;s�Z)�Y6�`��#���Z��mH�q:8���ܠ��^�ѷ�K��=w�E���gT����fCj�p���B6X��;�����:b�G4�}���F�`Ώ����q��`��
���E˝�{��Q&.A��N!��M�4h��m]�5�$υ� ����i��+φ䷚�Ë���Cr*U�v�?g����q&�Ъ;@�Gp!�΄��u� ��C-�@k��V�@� ��a2S��M�nF0����/��yD�Tq�[;v�\�V�F�]�Ҫ���(; ��⼛�r����cE>ʔ���5m9��A`Q��J@ t,�}���Z��r增�LZr��r� �}���l��9Hm�v�@���c�½mQ���T�<��rxzζmN;��]�.�U�sp�f�%iz[�u�Z�@8�g����~n��W������c�`���S9Z��VYfsØ�&H���}�p�8R�������֌e��q�$W>O��u������2��찑�5���J�IZ�=&Vh�V�V�K�d|r������Yo�����j���d��r��-��xx>t�`��N�"ѹ���氋R��&���u�;3Xp4ۮ+!}�ͷ*��E�fS���+�����|)���R�����'�p A��/D$�0Q3���P��0�8&�P�5iE���4I�0��4��D�D�m�AN�\�=������a��>K����v{rpp0�h?@ʷ�륵Zm��EJ�yX���������_��'��_�ԷZ���Η4?��|��V�m�B��)�x5�pI��zt�`��~��8�Q��pD;{�&l��WΨ�u^8[�w$�,}�XZ�S��9�Z�)��]�0������K�D�B�`���.5ipd���Ю"r�˅�p�� g�=*�X���D�9��SA�����ǣ�e������c$���C�d�$^(Bj�9R�8L��T��o�+Y���GmR��7偸��N��]�l���l.�"1
��,s��\����EZX��#U�fe߾j+�p��<�g�<A
��\��b!�κ�u���q���H9dѷC=�Ru�2��6]�|G Zl���;��1���6�<�z�*�n��S�;�n�v�F�v�����d���A�|F�[��C���B�"���I�>7�@\��dF4�`�?%�Ctl��^����m}��9Z�9�r-vĶ}�(Mp��s5e{ݺ��<�nF曌��zm����U�ƫ��H��1��RY��;�bL�jD����0�a�X~z���'�}��n-W�_ݾu+��ů�zw�r�6�O�O_��K�doyt�
Lf���F��x�����(6� �;�306ٹ���%q*4|��'�m�R5�z�Au�>Q��2�h��� F�N��ә�~����Tf�RĤ0����+!���i����^z�q���y���z�����Y�����4C��bt�/[�?�j��i�O�Z+�/��n>G�bH�3�ݎ�1���5�5����y��r�6M����ֱdN04�!��
�5g�i�����B]��B�y�B]�F�R}����U�+�-U���rEb,��U�*FD��P�#�������dB�~t��C�T�H�c�����Ȏ=�Pk��{t��Q_�,N �;�h~�K�:PRQ�`��"�!��d���t�AD� =�c.��!�k(?+6�D��}n؎\�T<V8:�\(/v\�Pd�t�����{���S�f�KˢJ���Px\�����j���%:|nH�W��q���ȥ}��n�9]�r���~]F���)��H���e[��AxP<Z1z�R���gf�x���k(�tV�`����>=K�>)7)�M%k�lI�h]JRG/�-LfO
*�a8�����\'��s�r�)Z?��e4|^�"Eկs��s���r�^%l>��Z��"���S��uNW��!
K�Z��7"�Lв����I�`	銿[������;{/�5^n4�QX�m�{�
rg����{����:���s�ɤd�Hk	�!�k�y+��gLy���mtڂJ>���� 8K{���@-2���ן=�@���s.�>9�Cz�¼�lcP��E��"��	ۄsF���>�m����?���;�5��F����w��m?e��"�ԟt���^�}�o���J�� ʌ~�K�ڄN�z�:>����~�|����҃�SF���m:��'iZ�Ҡም`f����Ȕ�p���2�3NK��&����u&�P�C����l�{ħ��h[���)QF�$�,�b�r�� PW�W��\���c����!�L��C���E/��''"�	o�����a��,�X�(�Ab��}i*�)S��r�!N�B�M-C��8d�<���f���pH�v�b�����2/ӌ��D!te�A���` U�sR�����h�γo�6/.�ې����k�V��s�V"s�z�/�4Bׄ��$K��U�wHx/p�LSe+�3z��.�L�18���I��3E�n���}��Z�i�8@��;7io�!�����9��%��|%uy9�(��|��%�����J�������:�}y���/v�i]?e���NO�:2��"��:���W^C~�:������o�3lI�=�(���.�&�� �u/���䬍���z�9�r��r�*-S�{�j�z�Hr�%�7��rĎ�9������_]l~��O@�s>�wo�������������ԇ3%�����5��0�X�g35��?؜2( 
J��oQ�o�qx�j*�Ra��溜�Ɇ�e#9[�s˶V�e�{�i��.f���:�56����V�^��>�4�����꠳��Y��;�yk�����_�^����{��n�NO
���jE��6�5�G�o��ҫ��!�;M�y���:;?�F�@�N��꥖�>UGj����vK��Hx�`X�PK3qR�4���B]s@���&k�d��Ć^�.c��N-���FB�-�:��9'G�����`�c�(��B�e4SJ�ES�\�oU��;�Z=?R��LwˬJ�x9(C�X��&���SR���m*oW2������s1�B>*e�u�
�j��é��U��Է��H�^8�P�U��)��HR���f��ھ�(s]��!m� ������I����R��>�k�gپ'���%72�f�F�e�Z���z`�O���n��>�W�`�Ǚ�7��(r� `O����!�y�޾�G�I�jH-ޓ�Ģ�����l�)�����������P*��
�?��-c;��38?�_��7�Og�맞��y͑G�ǳ$�I�mlx�25Q:��k�
��`Jj��\RX����<Y%�(�@SEF*�ˤ�r�&[�X�t1^I��t����R=D����w��]h��%�z����>]���^=�hr6���{������,����ò��c�z�=u�M�HR3��x*�2f�H�Փ6�D.�z�%�A��Y1-�ʈa2�����a�В�|F�a�s�L!�b��N�<;	��ҨZ���o�o�4�����bw��Ѫ���ᒞ����W��G����=����Qa���ޡ�?9����ZNΩ]u�w���G,�l4���zp�`g�Hvz"�L̓].f�8�uZ"�����3��U���,�h�l�(4#-2�����~���@f� k�p<��u+5Jy�����d�"�V�3
1�ӏ?�=� #Z�U�de��r8�4}v^-���6�"~�	F�Y�S�]��0��m�t2����Ʉ�qo[��Z�B�O�*� %u?�7�=~�gk�\�z�p.��bt$��Ò�-'I�
�H>7���8�Ę�+��H�ҟ��J2�5L�4��ɹ��i>��>�02�~?3W�����	�Y!q��[f'�[f\�YU�U�B&-e�X��^W�w�Z��B��U�++�DO����C�A�*ز�Ch�ͫu��iL���?�W^y�v\S���|�%����AOǢ\���U
櫵���{��vKͿf�W���tb��jת�G���R�WW�5'{�_�1o^�L�W�82T�r5����X.� ����FT���oR��2���f��w���18@�����K�%Kר8C*6�������_�7����(�s��|t�ú�N�uk�\�IZˢ��X��ʄu�Eq��ؖ1nl5T�|6$[;����bO�;xzz���3_�1r&l;b��bD�����=��&�z��i���q�����ӛ��;��9����ؙO�f��g��p���0;�[��*��&�����Z@����d��?��L�b�;�$�g�Dmv���um-MU������n���mh尵(���\�|��bO�ʕ�$�ZC�1P�a5�PR���YR�4��h��{���IC�ޠ���kt�p	?)� ��
�4��nb�6�9��Fᜦ ��q���[VU�#�峓p��G"�"�##K�K4
�l[��彸�K�P�V�9TZ��©�(�H6�XH[`gzz��7�)�\��VH�(J��*�]H+�:�&���]8Լ����N�#�~?].�]tw(��X�Ŭ�����{AV^fu�JH)x-�)r��!���!�$����R��Kj�{�2�m'�6��L�@7G�4#Va ��{���q�r�!	1CIVb���v1��$���g�@���v�D���Ѣ��:G�yV���U
wc]f3>ښs]{Х�|y��k^}8Z5
+��HQ�/#d������������R�w��l�n����6��Sa6�|��!?�GEC��W�kK�O�q,:�3b	�ʆ3���v�����/��4��mCö�ۮ}�Q��V�u�V�>�����z��|ooo��^2^��[���y�u�;����N}�A2�P-����Ξ� 3�@+�
	�t��V<��������x�.��=��;0e$�h�E��Iq�s�P]w��v۔�)��VIDK/�E���#���V�kudظ�ғ�S1�X�A��-�L�j6Z"���p��`�
�q&�TQ�E��q��
yF�P`Bm�H`n[�ۑ��l�x�F����vA��7l9��$�W,m6���b	��\�H��J�f�N7�,E*E/�x��{����1����ƺ�e��\%^�Sy��&�5�6_�t]��������U�u{�^�ޡ3�g	tR%1a�A�HaZFb�u&��LaS�����,�Q+,����}��O�h��H�ӳ%GL�ij�O�Un�5��s!�|���:ڍ������f{O�u�#Īҡ�_����Ǥˬe�e(M�"z�֭����������o�g9���D�����6�ڄ�;�qvRfC"�pO��u�"%|z>[ժ�!�}l��Q��:j4�?���~�Ѫ�w���Vc����������X��˧���^�_�/.V�S�+i�XN*�G�L��^=v>�Wj~�p8�ќ���b��Fk�Z1IJH]bo��G�3MU'�
���i/�y��C�0T�V�B^O1����)�!m9���5���X����R�ơU�2%4�LM�I�hC��Y��z@Z�@Hk���	�^�s@k�s������� /(�UR�4�ũ�ġ�^�f]�=W���!��R��V��L^�̵ӆB�8u[ى2�U�>��T5cI��MQg�F������f�:�����Ѳsb�s>��z�	�0�l����BDש��fr��v:_xl�Q��U=WM �}�Z�T9�2��� ��1
�:�s�:7��3G��O�v������Uщ��h�*K�lU�v�e���k^ܧ�g�Kܕ��$g]ڄep�[L��Rn8<�Qo�db�:�o�ş���̓���!mݼ��uDH>�tRbx-�>���Ԝ�	2 �)"}P���j���7n|w����j����no���Mذ�>�d��im��j��G�Ved��&��V	����ϩ�����6X�ф��9}�����]��k�2�DE�jR8�W��A��rE�:V�R��SZ�"T��uJQ;*�e`jAK�Ɛ,�����m�P�c�ۡ �kWs郭`�C�������'�)2$�x1�u]��ى�7������v���iz43�\O.k|.̙�2v�F�q�*}j(��D�U4�>糊|���R���.-8Ey�+}c���oFMЁ}��h��e�N���2����Ni[S�
jNJLB��,�9g[qio�s��eG�kW��u���˕��t'�L����T�p��J)/e�0�,��l�]a$�	����}G27K1�@��Ք"]�(%�ŉ�T��e�8ާ��~!G�$Nh�	_ �MG��j����$��;���՟��A��{�.����0/E��7Ϥ�X�	Z�H��\ mHst�z��7[���`��!s)u��T��)�}!b�/�d"(?x\5�\�o0���C�8����[���/����/����������-�N�OO'u���-~��vvn�v���Ǣl$s��ݦW�ަV[�jU�x�I�z%U�պJёD�Z� 7��98��È�P�H�H_��w!�j��fF�`���bCX�6;�~�A�Z���3�έ�{��MI�bt#D�"��ә�$��1���w+�l��p`z�	zʳU���(�LQ8�m�,C>��!j`�)Y�z\�/0e�xԵ^�nݴG���IՎE>ٴ�����W�0��HV�Ǻ��dP�j\5uݻ���{Z��������,�u�*�yl�e;��ss�Q(��Ga(��WW���R��Y}�ES���]��%�y�$�'4�p ����>qɌ Ñ�'(I��ixA�b�CN�G�~��r�![�7&����19�՚�@���v]���t�W.ұ�}�UҾ�/��J����T�_��IA�H�A���}���(�\�a;V C�O��U٠�A A�(2!B��|�
Qő�2��`|^z�r�в�����w�9�/��n����P����*Q�b�W^�E_y�y�ʁv-���"��)}С�l
|O.�F-ѭ��UM4t{
�`C�B�TrŞ�8�}�F�0M%5+��=ldcd���������o�L}F��##e䲜Q�:T�m	(#��>�`*U�	:�I&Д�4t����,���ٍ�o���^�a���,�Qn�Ѻ"C������2Ⱦ�|m��ǔB��n2� LՃ�v'5��Tm:�����E�Ῡ�����~Y�͵�rq�6\���﫦R;���}�rM���e��U���cH	vd�qq�L�R�����Ve?�V.ӕ0�i���t	 A��^�nHF"��aP�B7��ټ������jKS�s��/�~���x;;�d6�-L���_,�`���?��-�6�kY�(����k��Q���u��X�<$���J.��&�ש�ʹq�^����{F/���:�A3��R�j�b\.E��@�#��B��U��@���(�h9LW��ߦJ��0jno���<��������l}�W��N�G_y������h��'���S��7��m�f@C6nUQ����/��i�j�b���i��UhfcX�WNQ��\15ք#(��D9�R��1-�)�<���F#چ�v�}��]���K�T0������O��2�*A0)q1<��A�a�	���$[���M����@[Ř~U�@�F�Y��|B`d[��m(CII$]u�ZJ�P��%�Y�7��hKG���E܎E	Ҧ�\d"���Ē�lR.Z&�9���]�)��\L��#�;��ge�����j������Ȯ�ْp�Y�>��0+G�b�T�s��B�ԅ�nK<b��U������a֟�L��#����α*өnD�Ii=�Y|���#^KM�d�������|)�9���p�P���d7�ǺD�XWIee��nu1^<���o�\�g�Q�ܤ�@�x��!o����g��c�l�n��t~�v:F-g�c�S�]zprJ�^_�Q�i"��Q����������֛���~�w���?г��^�����t:\d�W��ʖ�w�MF���nt��_{��P��]����te�>5�-`��u�'�ơ0~Q�V�8�F���a)"pd�W�g��L&2��f�n^�=dT�@��mt�Ѭ�F0Q����0,����՗n���!E�!=��Qrv��0��e��C0��Jy��� �QS��sȋF	E�b��F{���uBG��Q��񫾴��5N�Ȃ�]����e@|1g�,!�U:�Tϭ-�Ut���Z��T����+�Ki�Bԝ�*�ϥ��p~����J&��BnU�.�����-�m���V��o�-�좸�$7�w1�(I���^��蒼�%�L�0O�u_)�)g�o{��n���X��S�7��:�+���N����tt>��_}�>|xJG����ݑ�1����yR��]�~Q�]oFa�O����B�����d��k
Â�6��Y�9���E�h�cߕ�.���'��-�aȄ��Ҏ�����7��K���u�Bo��̟�U��������d���r a{�>SC�F�6�_�b�V=�s������G����?c?%�J� ���I6����wz]QE��Q�0�d��QZ��ڢ#�jkKmGIF��@��e`IzY&NA����[�v*e�_����:Kd�e��G�:��"�T�ee�x�c�"ho'+J'�t���w�z�0�*u#��}��`�i'�>}px��QO�v�u�*�������dpN��]~/FB�O+���C��[�` ]FC��Db�s!e9���8��:U���4��6����Ia�ګ"_�kR���ĥ]*�Ԩ8�:����uCQ-FzJ&��@]�G�tp����*�V�����&(��Ƹq�#e��R���o� R��:�k���l����/�c�ܧ0L�6V	��"ڿy�������e��
�ѼW�˞����ɴ��MJюχ�6�7=��g�m�X%�1�3�*�j٦s5�q��y���Y���~��v�qhJUYU�(5�M��p����������_�+j�5j`(G黭5=��͎��/�D�GC��mUGAC<z-K7��r!��l�߹{�ſ���ӳ�Ԭ$��"Kg���^}�G�ݖ��;�dv�@�b��#���/{v�X�}p���4c���{�0��)�ʐv�h�43-.5��M=�G�,W2�P�*D��Qc"�Ԥ�������q�S]��.��N��`B��)�G�H�#\̥�
��[�c�Q$��聰�W�`_y�U>u* >�[�җ�P���2�4�k��A.h��Z)iiF��V����7 �gd�,�`'tњ�u��\[�$%U��m�~���JzU���8�hSQ�a%�(菟Yqu�J�!�H!#K�.s���|����"�/��:�z7V�*�
����BKNJ�E��u���"B]z�>6u<�����	iM�W�s>�v���S�dXBLg�;�{�E��.��:Ub�ƃ��q��Ss�S�U����T!���AȤ�8ئ��:�/�h��8
�p��P���~1Ѹ���77���֓��y��������F�cD+.(�<���?�:��#r+�T}���G!��t���Rog��CZ@���6��j)�
�aǶ�J����[7��7^y��׿��g�;O�r�8�m�d<��>&�Ќ��`�ڠ�AĎ.� �)�A�q�0���m�0��l�\�h�τ��-l_M�`�%MAiY:*B/7�m)�'&��PjEH���^q�8�	D���Q�-z�Q�W_�޸�K9#�t:���mgPQ�2�YR�Քke��3g�p2�
�A�d�Y�n�)-:6#Z>���7����]*	|=�F�<F�&��\FU.XՌl� �uBv�+v��
fHG��$:�״�lv$<JR��Y����O�䚯;�Z��`�J��2yb!�ʌ<K͑��eЎ��Qֲ���B�_����\S�E����`e����u��P�W��g�?��]7 )Dnhэ�>k�!�P|�3�L�UĎ�r�������ڛ_���?�R믶j�=z��j��[Xrzr9ﶱ�%6�'��/����E�{jY�'�e��7���uE��u��x�!<�^��Uެ?)�\���ب��}׶���r���p��|��?��6���}��;�f�Ԥo�-v� �������/B�uɄT��*���`���w^y��������)[�Y7^5�q��5�t��
�)��v�~��	M-���@&�i�E�����j�Ğ0�eʓ\[���B���<0-l�gF�j��JM�v�݉)U��9��cL�Ĉ}Ya�19i@����[oҖ������$�v�B�r�T��y���5;��|��Kv�i��g�i6�m]$���{[�������4
l����sT�dWf�2dX��͞[f��_ǯ0*�g��J֯(�JE����s�\��WhM2y�a�Q�v>���&|xT��T�^e��C6D�U�Q�-N_(d�aB�:�2=��-�5�X���g�[�@Z2x��l�heD�i?/;�͵i��Q�w.�w	H�L
$[�c~5����E��Q�O #��>~xL�~�_���Dj���`p�K�X�����\�~��=�c�e��a��������;Z�x)>�&y߶�e����
(�Q���J�������i��uͣ(�;:�h�
����R\�#����x��ٌZ�6m����1�f���q�
�G���:�8�2$��m%|a�������	=[O�z���a���'�0M�J��]A�H~rx�H0��5Ҫ	O���1����Qa iZ�d��q����|Y�2�\n\/�}�[���&� &@ٿ�e��oq`����P0���6�T�R��ӥxxL1#���G/��8v�f�&l8?i�\Ѓ�� eX��n7�ݩ������6%�K\銖y��m��� u�B�8�:^h>ǉ!�e�P�Q�p5���
��|d����B�\�|��l�[�� Mm�SuT�t�1��zPI9���i5�񙅣��!=
G�Ij��:U�*=�m$�]�i?�df���CkBWYs��\%4��sQ\��]�P��U�I�;�7.lrY7)M����m0�a�݌��ۢw��!�z�k�ݙT���̈́d'�Ӥj�~S��$�|uIA3���ٳy��]��1Cz�S�;|Ό���6<��_�����xc�\}�%�]\��������`��JZ<K�
�����m�&�a�
�;�N��?M:��X1�����`��6u����N����}��o}�[z��ƕ��(��<���3��8�&�f+������SF�UQC3e`{FI����$m(�a���
�糓F[j� �2/V<'�Ӫ����e����B4�3MH[��t3#F��jN{�Io޾C{�:~@.��-��26��ܒ>J�Ժ����x0"���j8�k�*�h�ׅ�D��mQdh���k$�Նquy&��h�DYYM��d
�a���s�BY2[w0�%��s�lqۚ�\�z�Ũ�e2����)�T���z]!)�4\�l�c@;��-s=r�ѸB�J�|D"ُ�JU$�5�.��ٸʧ���CM����E���U"�M"�t_�[�.���Ǯ?�^�Z���wK��k�0�F�R�C�Q��4��d�9G�Ԧ�t�D)��
ˣ����އ�{p ���%�K�?���e�"�m��x���;�f*NO���8�(�VDΡiZ��<�T���:���K�%~��m4=_��:T��1�z��jh��,@z�L��G+�O��5�B7����_�����)�*
��T|ŐD�7����|D9�I��jUH'��m�L���pg�o�޽{j�c9���j����M�ه�GS�o%��َ��l�>�j�G��̂E��d�ʌaX0��
ZU�Z��8��@e��)g��%R̐I���PKC�Z�"�T喙=���P,����n��?�ƛT/"��N��"��F��_�٤���H P�� ��|2M��3q�Pv��ۣ�?��4�:#P\�HiOc�V���ޗ~�D��v���2�'5lI�f	^� E8m�!�k)�.R������J���(4'��2�"����q�} ����l�6���;�N��L��j>�<GF
���)h������+a��ݠJ�G��J���he��7�[�
*�w�F�#����XN��:���~�I���)KR��!�&F�X���Bw3J�#F��n&���b�{�������tdOv�=*[8QR���z㍯�G}D��ݤ�b"��y_�&��2���TD+r�G���D/
W�l!����ɇ�t�h:�����-q�I��g9�T�gZ���:P��H��G��uM���Ys�7�H��#ԆV3R�]�8d�P}A�a�ْy��L)&�WL���<�::=:��Zl|�Y�΍}z���?���2��	#>O�b�O���/����{�ޘ���v�y�4\�4�8�~�K��&�m�b�0���ڣ�2�i8����H��,Q��h���� �Q�GKvFh+�Q��C�N�Γ���Q�%���ma�g�1��1�yA�
B�gJOjJUG��8/�Ĺ��M�m�^�٣����Ɋ�������6�T٪ќ�2�3�ب���P�P�?g�ץF�`���-C;���pB���R�Qǋ��,a�l�idf��F4�aM��qL҃k�CN�ֹ�?3$è!3vk���o7hp�Ϗ�Qt��휝�ɧ���>��c�D���A�ϟcĎ��s@��[�\k	��FG�i�ȿ�N��i�y��!;����z��A�RG֓��`',ȋ�=j�T�T!N�A8)sx��Q���)�mO�z�v��sp_�7�mS�rq?��%�mH-  �nh:K���C"�Uv��p�}?��S	�������w@����j�s�I����/��/S4Oh�U��ɂB��5���X��>|\����t%��3:Y��yj��(�x�C�1������s�\?I���d��x-o�'�:�4j���V?�M���$�p�G���������)�L(��=�1��/�F��!�=�ʋ�p.hΛ4���#R�]�c*����֏v��Ϙ�O�rR76�`�!��uٲ�U|i�Y�����y��%h�V=��M�QHXR�1�2˖��ؒo�M2M���#��g�����c�I�x�D�*�Ҡ�/��^��rg���!�}D`�ܳ�Q���7�͗Tm6��xH+�Γ(� �̤�e:Ju:46��q=�d���g��)Gm�P䙂.�a�x�R�s�ɉ
��2Ծ4]��eS��FR�ȨV+��)��zk�h���|(�|�s$L�gt�1���&4_����Q�J���1���B��d[�b'�9Òm��9�����i{@�*�%�n)�ңl��&5LD�|7�N햢9p�H)��%u˷'Z�'ݰ�����Ig+K�r.�Z�0.�G�W�!"|��Gi�\gUV�g!H�����O�͗���"CU��ùı�r���'�"�D�{}�7m����3q��a���x��ֹiZ���"}�
&���<�B���ID-�RܑnQz�*�R�@�>2"��xp���e�;Z������l���F��R, ���76�"�8*���N�����w�����l=իR)r'4W1{3�;@�2vF���b�VrZE
Sُhk1/MwQ���+���v�2u�=����zg�Al�ؑ��,Ҩ�"*a����h�ªG��j����}��|��Ɵ�PX�Nݧ�xN;���>�3X-ɫ����0���M�hĎ	ue�P昡��bX}Lm����RȨ7,l�y�nX�l��.��Jd#/ў����u���h6��G�>�=�OМ��<�%m�`�?�/d~���Ph��m~�hI�bE7�]r�5 �-C�հr��T�Fi:��v�A{F�+<0(W���8�%�}T��Ё�՚l�S:�⚁7�vvs�����mq����`��S֍��Fl(i	n\�&�gE�����?�����åz�I�UB��чdH
3�,��~��F����do8z�e���[�������b��42M��_%���>�'���M��<�����+��p��(fA��=�P�p9?���n��R�Z4�,1|~��ާ�����S�ߧ�t,�QՊGKޜ��9;׊"4��h}G�3V��v���;����7�l=ի�^.#6�K�h��N�)2�	���P�6��
J)I-j�"fy��*d'dH�!c��q�ݎ�j*�TDԮ;�G
N]~|n+�al󬐩;�����^���Wo����ttzBm���+U5K��X�+FO�d4^�t�����HnﴚP��j!m=h1J���)1����eI��v�5[22��v�l;��/�kن�Z1�Q��/��gi!��.�s>-�F�����j����V$E[�3�{;�O��"b���OSR�('aFW*#]5��R��_�J��֨KϯY���V�f�K�X��l�բe�B�Ņ���:׿-�y�Q^���ق�,��L_�����Ij�|d��!mU�tcg�v�]>l@}�b#��L�Ǚ���.�k�v!��\�5����Ř�?��g�h������xd��ٹ��n���}�j=������':jy��Y��c��a��K�u�
 DFn�y+}ʗ�4��=�0�(�V�
:�Je�'��w�!�/�~�/u�p�67��p�Y�_�?�je�����^�wN��S�x?fn�4E�	���5�`���tB���ڂQ;��e�ju'c-^�~RE Q
E������j'7	E�vhE������9�ޘ�Sd��JF�ttN}3�z�6ݮ?�G�xE->��dJU>���n�x��{0�;��O��p<&�֠hOZ.��yZ�n�F�h��H��N�B��ūS���ٙ�fh\�B(mK���M)3"�ʕ�u����XRg�u�z&�m���9��v]�W�|�6m1�R�,T ���#�f7j� x��V�b߇��
RHE�IZ������ً�b��b�Z=�*(?C^��K?����Y����� h$��o�@�8{�C�T�(�LQNp����k/>G�ݼ�`c��G|"�2A^u�%4�l-"8�Nl�͊♣}����ll�ٻ�i��&����o~����_���oΖ��y1#����\��F�v��)G����+Lc`eF�eE�f1`_;�ԙX�b�����d:��'/�e�=��#��{?��f�꾚J")RlQ��3�0\_���bk����Tjg[�Χ����g�a�̓��2L��S�:l����'����R�d�rp��qeĝ��A�1�>�T��Cz.cC�v�1;�Dlc�(�F_�qyDc̗w�֍6՗C�B}v���lIy�"HӨ\��#�&47l:�/�[����~VKIcW\O�p��� =qaVh����p`Z��3K���Rǅ��:����Vw1hm�f�F�傑iB�����s~���W�0���ft��M5��� �/�?C�j]�B��9��1u�=q�QΞnv�<6�B�Zo�B	��ϣԒ������ 7k�8��[Z����Z������t�tS�jFpmsI	jt�s�x?8<����{�ַ~W�s��Ć%���3D�Y��R���ԯg�g?�N�gJ���ܴ�#ۈ�:�b��J������s����1��"��C��o��#�W�AW��׊7�ߏ��+��?n·��Se��.�$���Vqq�}¯�->������_���âG�O�N���kVP���D�@�Y����.��JM.�J�J�*�����������}�g��`My�۶�؉�I̗�����t6�0�h��8(��@�P����FV�\&�5Τ�QO֤�BT�,#Q�y�z[J�O.m�0]�w�箺FJL腭:����h�Qmz���1���&sAm�WeW�������Z�Ci��w>��2�J�%��⣀��:�n��F��`��u6�e�4,lq����kA���HO��s=[,7�S���9GJ�����[`@C�B�ytT�K9��WuXi��s�C�[�'T��0H������G48?�����^o[�2�O-b�5~�Bq[�K�o:���3�n$�)d"LE.�6��������u+���H�gC\Hγ&���Y���K��r�r�HO`�h���?��h:�9[�	5�����L2*ՠ!ψA���I���)^?SG�������|J�m��|�[����(T��j�z���q��H���ڼ!z������f�3��0��b��9���*;1:q�Jř��S�rWIbG�Da����N�9>V����ߜ����>::�w�w��j���Bg>�����)!ն�͉�H���^!8�&�������}����P��k!�3�K���S�D�a� �
��(�"A�\*��4�RZX�0�<�&G�#xM�p��R��\�D��cQ�m���Y���mz�F���}Z�#?\���o����Y���������rA��ӌ��xB{�f1��tp&{�~S���Mh����j�g���'�Y�WPT�f��Z��t"�
�����Z�ȉ��8MՏ:�㹱�+i��p�u*��E��)vL	Jex�-�i���$��	�E���I<�f�Zk|���O���z�.���y�yZF�|xr���:�+Lc�Z66��T����R�=��7��:�	�Ua��v��o��mؖ�����j�S�Ւ �16��z��m1և�2!�������ҫ��'�d��fD����[�Ԯ�����Ϋ���y�{����&~���
����M?ڔ�,0��1^KG���������B�� Mv�ł���Z�G�U,�̊�Ԏ}?cd˗B�dp������xt~�z�w~'~����_��t{�5�t����ww�ø�4�~�Y�h 	9��H����"��4=����S��_�=�IV��&9;7�C=I�B� u��cI�rƌ���T��&e��pZ� +�ٱ�tP߅�#�~�h1���$�a�M�BӐs�.�'X��Y�T��]���j���]����Qی)<}H�jF;�%A,�s�)&��gqL0����rJG�5�U��7���`���D��d��ץ�y;���L���fr=!Ɛzg��K��KH׺N�r�<�s8?�7�v�?[�2��h���%y59ҁ��>;��D)�AF�Ʉ^|�v�Cjz&?~E��R�#�,�4���a1S�����N�邾��`86����.�1[:G�z�^�� 6C	P�b,����jF���/[;gQ����&�[����jF`�>Z�j�fD�[����$q�$��VP�T|�}�(�d�Ѧ�jN�ɀ�E���6a��R�rI�JD�N2"�dY̼R��qL{L_L���x���8n޼����/�0���C˰;��49���nb_��t���m����-a�����k�5m�M&��r����2��j�q�n��
���-�w�Y�~�G|AOy��-Wu�B%Y���ܘ�9L_��FKG�jֆ�V��kY��/�2�z���_y.��R�Ø1��@$��	B	�\�i�u-N�,s=���l�Ȥdkh�!�HK	#^K1�#�N"N H;Z���t���_g'�|å��{TY-��: ��/j����
�=#���N���4
Cr�5�kJ�0ƜX~Ϫ� �4��ȩmQn7ة�(3}>6F���$	�4d��&r%za]�Aj�����##+}v���A�Nn�d��b.i���=:=���!�}�����ə�V���9���d�B�S8�	2�sS�Al���}���XRӧÉ �ę��''P�$���"��̭bm��?���G���>����$>m��E��������~CՑM	�g�0u�2|Gfl�EB3�4��C4�UI��!u�wB&=� ��7��jPM�ɳ���dmmm��KG�љ�N��ӌ��,L#4���-|��5`P�f��j_�Y»>�����o�?��f3h��'Cϝƌ�ϵ1/ԍ"ՋK�����4A�VVb��cnZ�;�G�_P����,8�$K�y�K�NZs�`���v��A��S��A���LOv1�=ߛ�%!���[�n���N�A���u�&��)����K���ӣ���L�\��gG����i�^���!�Z">���O�~ď=^��6���"�[��3�beV�f�hU�T(a'��� ��#� �Lƚ�Q�Rlfs��7:[R��/���E�,���,O��V���i��n_c����3>/$����	�>?~H�Z�v��qS2�PΎD042�_�ׄL�R��zݣ��FN;r<}����е^�U��	�̦j�*�5�E���A��3�/�h�Jֱq��p���U�'��Z+��h�	Z�;�s�r���������@JJ���Y��͍6=��L_R�̧G��� �|�3���h�dQ���#�R�l
ǞAo�p��@�,d�s��j�Y���Ԡ~qV!+˴�yئ8Y%���E�
d(���@Q�T�R��P�H�IZ����Cا�0jP�ָ5��mR�fzo�m銬՘�񐑬I/u��[m2N?��lD��`���D[�:E���.;F��2����Nة����|�	�,��EP	�_�����8SW�T��a��j�*� S!��
X�������GM"2�b�Q�	�k��3�[�J�"Vs�����ծS����OD�c{�&ջv�U	h�����j����S��������z��[�J��	W|�*xcZR��ȫ���1l5PH#[d,���r�h�*�a�ed{���8Z�����'��˂��u�w�_���ˣ��e(ֱ��V?�K68��16�΂���L�:�2�,�4a�|7��P�g����������2Ir̟�b~��N`<!���jA �����q0�1�n�7�V�=[�0k�
�>�p#-�/�l�5�V���%�S5�Q@����Qgq�`��]��O�n��2c��C�@(���	�d���s"��N�~�f���Z4|���8�Y��*N��m��Ă�������و>=��t�j4(cg�X-�o�r��N�����<��%2�C[�����Y�R-'�^J]*R��9-.�܋�g���3�ѿ�����t:��0�}FھL���b��
�M.җ���!�i;J�PHH`�����Z�l��̵|A�?g���m��S�koI�P!�������lE��Xk������m|ׅF�k�{�֎�q�I�Wu�v�����t�dc�x��q��
��F�&��J�V���֢,����Sz��������g��'Y�ڲ�n�f��H
j�+�U��rD�<�Ƈ��7�N뢑^i�%�No�	_��/�jfY>`p�f�IC��=�T"��$�,[�mB� �K.�>W���Z�6�eMO���Q��0�Z�).�j�H�^!��8��/[Rێ�nӥ�ި�[�P5��^�$��,����F�N�,�҃pB�gC�rB� "w�)�A��fd��=aZ��dN��%�:���N�*�6�6|���R�i��[X���Y�Mf�fZ��GE�p�@��x2�d嚢���Bb��s�\�1F^.泵�f�JV�c!�!ԯDA�N���9`�ΣX���,��1�k�����2�T�,;�Tg���
mG	h<�ִ���q�����qu�ϳ�͸��.�5��Ǘ߃���b��l�ҡr���Pë�6E�IȾ"Ү�LE�ϑ���Z������IV��vv���y�D{�`�e,C�6"��Ck_��el�`���&��(�l�g�fA��2|�Y��	�"�
Z����	F[��E���>���ιc@:B^+W�m
�[	/R����|���نt���{5z�mQ/�P>9�.�?z>1@���[k�
�F��CF$��h8���S���6�dr �1b�+�5�)Ԛ]>��n���F�Y���n�t1zWQ��3�I�	z��S�L��3K���'J�s�t-U�V<D[f���?Yǯz�|J��;�#)wC�yL�/r�=�Y_�
)�jC�öoK]9�Q<.0D!�ϗswa�-������<��!��J���̄d6li��j��H��z���u-9�'ޛTV&.�h��KR����q����452��!��t!d �1&��{d)�i��˒�8�	6�ͤ�L�>-v�|*�g����5����V�	�P��$��y���w�M�j����)˶�j�:�s���L�֣k��`�ؚlQq!�8E_ͨ��T�!�`a"zh1UFt��Ƣ�EU�rQuB�?P�mJ�T���h��zQ��1����xJ]#�;-�^�U���|H; �c������-��ޠ(��䐚M޿���޳I��:<׻�Y޴�'@P�Dqd#�ڕ��F����F쇍�_2�_vv��B�1�f$rI�PCR�"A�эF��.��>�z���ެl��Dt�^�XUٕ�7o�|���<#do���p:����$l>�B2 ���E�Q*���t�>H�E�d�La�`?:��"�K���4z�M_Đ�T�C�������J"� �EWxV'�,�AB �����-V��ıv� � ��m	d16C޺��u.�,b!��VF
\�����y��j����<�i��Z��o�֛tH�m+�"�Z+=Fi~.�trٕ��f����t�˩!�X�������j��]�������$��f +�G"e3�DJ��3�1���3-��MPqJT���Pf�o�@|]]�u��e�9���C�Ի�x��kueJ:��ɣr�:'SP�~f�? W+��k�`�G�:M�z��:Z�p?�.�I�&)n�����1����G�DF51i8U��K��LDM��إ�����
��5��NI[�$t���fe-�a\��AX
��ۃe#�G�ߟY�ᤎl�p��]�}������6;�xPj�Kf�f.\=�؛��-�@Cⵝ�dX`򜸉��ϕ�q�$�V� �pE��&�,�! �m��,Y�G�d3'��h��8y�-OdQ��O2�qK�%���R�9� H��"��c$4c�D,���*��|=o������,o�a{wF�>���)�'?��F�ݝ} ��샏�)�$.�`�s�x��$�źà+����h�y�\��1r�^W&,)�.l4��gE��qmT�o-����Ι�ʳY�0+PIw~�b6����m��s|�� �&<��Jn��aΪp���EB?�I�����d��9䕥�0wẎ�� �k��>H��v��Q�aO�]?��̊�ֱ����s��/M����k%�&G���C�:��Lq�lY��C'����a�Y�NH{������x}�m�9ON�[	��Pٖ"{("�Y���I���������Ru�*�e�k�<���&�U��$���}��1���[���X3�q����6�í�(��{>i  1	��C<Ɲ�\�O`A�E0�( �͓F}���z]�y�.�V��!M�0N���}���r�/A�ʬP*T����#0Eg*1��V8b�e�eƼ$ѪC���2i>Y��?���c��:2����	���K<�B�Ԫ!�RZM�b�#SD�	�h��fL���IZ�	u�{�>�GQ1�w�;�Q%qR���	���n͚�:d�ߙ��^G�J�}Ϗ����L�`�^����Hi�����,j6��OH>�0�f0ӵ4� N��$�����g/�#g�����]9����z�o7�,;�]Q��`MD՜:�}����3����@��$�H�s��`[���~�VΣ��<=+��p��ts�f{7"�'����R��f`m%��@�TI�o�!w����E��1��d!8y KZ
�U>sr	6�e�d�Z���ƅ��<s��R2�N�1>v���K��rȞ+� #��d$�X��m��<	�� L�8�Ht<<���DT(s�n��h�J�b��M���+ˋtyR�=^)L/��KVV�񈓪S��R�t�DT�}��t�
�s���z�f�ؕ�H�N�<!Z�_Q����KG���&�Usī�ʔo>�p>��e�^�[\�iшU�����@b9�&7�l:x��1оוہYo\W,c/�V�a�,��"��|J�D������� N{YEd�uM=>矬��aZHf���CSٮ�U��i�D{#��U)C��vT���9ˣA�,� ȸH'9�kПN؉�F�]�d8�_��<�q���#�m]�:�F��m5�B��X,=I8";팆���V�}�:���G�Q�oI���n@Y1I�=���r}���
�:�� �	6JyaȞ	�F��ڼ��l��nڲX�<�̽M9����R�ө��4�4�ȃ7oB8�#	ܫ�1�u$s'-~�I���)LQ�	/� S� $�K�YFӟ���DCo�@����b��49�*����V3� .��]���4���x^bYdd�[�2�N��ΐ�n&�xg��Yr��M@�7����,����V���ြItb�4�C��r������y����k��hI�:�A����<^w]�³8�g�ٍ��X�KM���y�� )!-۔z�q�h�"Q{U�%���,Rqx���
�- ��6���:<Z�੦	i!����[���]b��ς�c�s�';���3��}�׶n�X�!��,:>"���"I�Bɽ�}Ȑɒ�wu�$l�S���!֚x���c�XZ2ϊ4q.@��΋���yF(''nN�hs.�<8�Bz$U(��M ���%�����S���FS����������%�u3��f<�4� �u=6.OrQ3�3>�w8��cB�i!�o�Z�	szi�P�}���X�\)@�fj]�5N�j�=�-|wܷ�N�Y&�y�exp��h��y$��ݞ^s�C��b�ק��h��*��a��������&,�긙N�Л.�UrN;���Ĭ<�vQB�[7V�A��%�7^�w%֪00�w��4X�k���8�LF�Z�e�*�Y9):������\xb�O6tx�.�3>���MX�?���Θ���ښ(u #!������o�Gp�������m����"� ���N���N@�"T8�`-��~���{��-S�bL�X�"D�7d�oM#�����ϖ�4��-~��>cI�*G�p����C���X_Z�@�¶v��%O�";��+ի	@&Ȅ��:h�X���N��1aKC���܃�d	��م���Po�t#ɹ��+��`�������+Q��ŎJ��B*��vwc<���E�~Jyq(b����V� 2x`S��@�>�RY���֫`�z�IN#�QD���� �J�t�������_~I���f�����K��z��UѮ$?*�͚{hS��1>I3�0��N<�|D�Jh�B�x�$̄�v���C�Sh�'�e`��S�&�62h�#�{�#��l[x~�lTg��x�N����Cx����L�+����=5��V����
���[m,�4�a+`/��P��d�~���w�*L�At���
e�9I>��� �Hz�ج�9�`�����^(m�H���s��m��Gl�@R���L���Pp���/<���=�LՀ�B�3��%�"N�W�Z5QϝNf���c�Ѝxt	r��:Գ's����ޒ��m��bČ���|��Q�<�u��K��@�~Veqqj6���Ms?̳�v4���z=p\j�iA8 (��ן{���d:v�0X�ͅ��c��O��N��������R�d
�GZ�J&F/�����ܕ���J�&92�Bh��%���,vY���Jǰ����m��C�����`X6L�cd�>�<za�x;�ׁK�=p�x'd��蟄,,���j�fJݵ� F��q
��'Ā�݆i�㱒:�`�2��\@7
�+�6��K��|e��+����퐩��k�G�
w��"`L85�ļZw؅�h��,��)eL����+��j��\����`�GS�H�̨��cV�i���Xw����0�Ge�t6;�2�z���h95\4@)�Ƴ�+Kud�\|���2���&Α�߅�{X�@�~��_=q�F|�����3�����uVV��]H{}X]^�2�x<�J�
�;��y������p�>1˲�ȉ�{/I���3�p�x:f��7f7V���	����L�p��jM0�E44���?�B��jJ��Sx�l��L1��= t����ȩPC7a<�yA�f��L������Lv #C%fM�R��3���Uh"���X{c&�T{}`�X����k��Ǭ [�l�ŒhH¬�t��Y;P�6.;�n
�`��#�y�-=\��'+���֌ٲ��yvӏBN��z�!��1�y��X^f]^��ާ���,����4�C�\ ~���,��]߇?�2�O�c�:V�R���(S>�,��*l�I�m�Lt�n�����ݮ U>���wN=�^P���a���z(#a෻�����ʩba"��p���[�� +��yr�ۂu��X�R�?�񨵲��������"uf��l�>`d9f#�M�"��~�O���=���\K��
��'fQ�-��S`_4��&+j"�:���]�T�ŭ(�
'��dɿV�|0qs��)~�aYO�L͂�[6<bK�MAB<8�x2bPh�Z�L�$)�q�<�f;�:^ ~ ]��u�U�4�ㆪ#3�ܣ)Ls�����@�Vq�$�}��}J%#1���&8��R�\�͏ff��¬���V6{����.�SRJ`��3���n�m$@�` Bƍf��~�V`����)�����q,����I#U�
T�=�t�Ȗ�>�k ��\t�|�+��w�};��;L
�f���v\�⬰<s�/z�Iz�:�'Ӑ��]�H�1�6<��h��r66ƫ��wiw��m��1r=�̧�Mb߃`4�%��������M��_���Ž��������k����������&�B/M�FK
Fr�r��ц��V��Ud�z8�f.,�9<�`���m8�{zcڅ��&��J�s׫SmB�Ն0B��t� ��t�����؅�j�&�d(K&:�-ۂe�D�`B�͒j���S�x$��*�ꭤ��(�ftguU1'���~-��ł�E���tH�y�eL3�,Kx�s:��}����Y�N��l�Bs���*���Hic���疬�z�	�Sa� L�s�����t�"H�܇�&�U�� ����<Nrf�^��c��rN�w����k����m������,��WY mi� �&H:(%B>��]�eVbv�u�p�u�n[�ښ���;���d�љ���K��Xn��x̛��ו_��=��y�����Ϝ;w��׃����v{�[671�3��DC��/�F�:�Nc��I4u�;ra�҂5C��6O�R�A��!1�.H�1�q�C��ˮ"(�WL�=v����)l�F�f�o���d0�a��#�1���$�� 3��8B$u�d#J�5H���JB�BP� x��Y��0�!2�MDwP�,诖l�����1h�R�dKW��WÜw��@�ܐ�3)�#6 
K�9���7�-..2H�N�G��g<u9�L�QA�R�4�S6���R�WdNS�{g�Q ��%6*�-)�;A��џ��Z��T`�f�n���;���v������?�H��d'�U���3џ�u�`Y��}��7w^�Y0�eM���t
~v�$\~؁���K9!��a�V]�vs�������J���Fq�K�,73E��!�˖��u#��[	)�����\u���^o^��! 7��@�Y5�rI7�h҃��.��*��z�d����S`J�<<�x��\.��Õ�z��倄�-9�������#cC�H0r#`Ne\�>>6 ���06�%���2�e��� ���.b��E �jQ�6K9���	 o�l���6f��g<gͶJ1w?��uqcĐ��(b�
��)��Ʃ� ��F�7�w^�jOd�N�P,(�F�~�{�h~�I۹�K�L���!��5/�\3aMǂ��^z����w��!�Q�L�X����4$���8n��jx��1�~�%-=1�񣷆ۻ/�����g&��Muơ��7�Z^��K��Xߨ=���k���S��|��z��?'��s?!ʧ)���g�0�K��I�0�X�B�s�i��X�tx���I+��t �7��u!<��j��{	���K�\21�L' ��|Q�}sw.��p#h ��>����N��`Td�S?�2Vϰ��+��T�EV�_$E�FoH�G%��(�*��Y�J�
w��G�����t�?o�2�v��l�^}���@��L�Dƀ JD3�*�J�iZ�Z�/EO��քl#���2י��g�Ur�!�[�1gU��U_X�F*|u�O��K�Ѭ{9G��v���>�����G�B)����
�Bb�c�H0y��������f����W1b~l���6+զ\�!�ɠ���m�!��nWYl��ݩ�O�n�xA�x�Ep��%2Ǣ\G����;c��q��<[MRĜ4%�����DPW�h�b-�i-�u5��ہpgb������C�J����xĨh��f?{��v�
��{��&J��Z&������LL��$L$%$��ZO��Ģl�$mT�S�SR�3O�g,������+W�i��U�y���7GQ���ͽmc��-��h��$��cSz�w�0>�p�aO�vxq����U7��Q�������ڀ��m�f����(th�kV&qS��0%&�}K�I��ґ���{V���~���Xhݭ6{�c�]�$�I�Pt.%I̅g�nf��wCF+��Մt�\�榟ooo���rx�9gתN:�u��[�س�c@i���|�y���ʙ��t��>�V�t�a:p��%I��ʒ�h+�3f���h����p4�B�E��Hcp�	ٟ?�d�'* W�����݂*��!�A�Ch�9�&�G�������A���V�vv�&P[ .@ѿXF6!c����Ff�&w�.�nµ�}��ʐZ-H�6���X^E� �QȀ�r��̚��=�Szb֣��E�[��:bis.;��51�C*X�8�R�X���1���`���iZ��#���%I�n�gR1R,~,���R�aaņ��m8s�����gBB_�� aS7x����������������0g PVd9�
��ޒ��q����~mI���o��s�;�w�j�\�"����b�a�{Wsla�^t�Ks�E��3�}��1�~k}}���?�;<xq����e�\m-����Աc�8���&�t*�K��x|w��N���@�J=8^�
���J�K
����:ePUIGW��b��@��j
���`�h�>��U8� l"?���2v!q'`Q=��c���#�Xh7ayy���A2������`o�E���>ĎP�� �94���a��-n�ͥ5�x)D�k?T��M�ZС����IA`��s��/����*7��`؎���ד2*)"�:���� )����β��N?�q[���¨ 
l%�����~N]�du�LL2�߽	���p��s��9���)S�Q�v��l4��O=�`ك�[Wp���/��AVؼA� �~'u,j��'��BJӮ�I���K�bt���
�Y�ѐ�۟�ڲ#`&Ayt&n]$[r�ѝ�6����J%��3�9�s���n�{:�y�!FX�*�r	\����!+��p�ܙ��J��+����������/�4?�xp�ܹ�Ңp3:8��Eu��9�p���(����L�ݐU���^~�9��g�]��bIj��x=xKUC�]Lm���T ^�� Uqc��'7$+@��by�U�y}h�=��	��>��x�)�C
>>�����
�i90�\����)2K���߸	}|�7�� 2p��Ue7�J����vYZFc�j<��j�!ەrRd�QF�Ţ�I��+gG5ڄ ����(����T)�Hs��)�G�����%�@zgu�l�
�s����I���s`�`��0�g��~��bѴ��U0� �; ���2�����V(O�<������!�����<جhv��[v~��^g[?�u��W�,xB���T��Vu`�f@��@;���sA{!��H��g�!���T�5\9�iI��&�ի�$��u/\�ݧl�Q#�-\�1�v(��j Q�	�������`��p���������z�����#� OSڨu'2ܦ:��l)5)E���ǰ�LɒS��)� �|Ē y �d�� r
�ά�d v(=��PEP�h ������1#d����o��0�፽=�LB�mB�j��R�F���P���s�R��b���Cp�:���@���R�8��"�əEnv�cR�d�,;J�f��('��P$*�J���D`�������������HO
J�R������Q����8 p�L]�8e`ee�R�9`���s*We�e)��S��r��u����1�3YBr��M�����*%�7�,�%����+i�3��u/����¤�n���n����	J���4�n2����N�e�r�w��Ha����?C�{	*�㱟hI�X��R�Q�[��C�G
n:] �!hI�@�&P�t��}���mv�A�
1� ����:xQ�Bidz~�`zy��X.w�#�z�n��Gvo�
11;t��:��!�nDֻ3�����@J�V�Y���~I�Z,MJ��$���ҕ�Դ�D!3Z�"	)JJ��5��`��6�u�ۧoYϘ�'!��3�Lawo�u����A�	�2�ఇ�U�&���.�AM�Yɢ��ϥ���ɏI�ý���}�8.z�H��U��N)� Yn��Q�$�ZQ�?Ze�EK��t�@�!.�x������'�� %�[����$�i�0���� #o

u�ha,��T�������K�ɓ���O�?l��n�cYV�L=5��D⺔Rl��	ٔxL|�<��!�2�k��.T�U�}P�	d�� �t1mhԐCC@20C�a8Cn[�#��va�������nnt���U��Sz�r�Sc��J��z7D*4o�����dCk�,�Dj��#��X��DXr�5�Ǔ��f3�-�� n��R�TF�� ڐ˔1o��Hȇ�-K@@]�$�O!�na�1A���vn��~Z5�x~�-�F�~�TW ��R0nu����ge��m*V��D��<�d�;���-�Q.*;p�8��x�ֱ�Z�q\���I1�U,
�T��fd�2���y�3��u�K:wn���_YO�?O�����ϩY��r̛	�y*T�~�+#nR���p��Yw80����L����mIZ��x��K�d%��Jj�I��Ҙ��GPG��x��t�}0�	��0쳔"�߫I²��R��(�FF�~W+6�2����v{ps8�d����}�!D&��6"�4�WxHGV����)��d
AB5�Bd���>�	�R��l�8]�S7���f�"0�J�WPgE'm��fq	OJQ���	�Ln�)dK�-�̣�mV� �+�rn��.?���4.U��I�a|��x�Ā�^����a:`9��m!��'���X���Ky1�"��~�۾����5�_����F��-��Ypr��}th<�KE�����m��;�pژ�1�~ky��L��z&��KIR�;�O�N���m��'`��)�§��M13Mh,魩;���_��N��s��^��!X_HlIr�����d��TͳQ)g�]b�2����~�����Q2u��7B��fu��aAn�S�&.R:�!@J�;�1\<8�+�>\�뀇[Y�;X@̋�s�n������C����J*G0
spc������p��D@W9M*%��fD)�%) e�_�b|�+��5V|�%��Ͷ���]Q���Ӗkf4��KL~�(g7���cJC�%�Is�Zf��j�(@��n�8h��,IV�t#���d�G*�Ѧ<�"�梏���p�v������DI83����戣4 �?
��0�~�������Y�+�ٌ)͏��z����z��z��WƣS�y^�D�9�dqJ��!��ϩ8�ג�ux�Q�Qk�֓�K����]��k���?�O��ޛ���>�+���,�22(YK���|0�d�
do]��`"�l�ר� ������`I""!�ҭ
�_b�4"��:�R�f��;�\�l'�6G���T����FXC��q#\�.�f���
�{]v�1���[V�4 ���16�T�S�j<SJ�\�!������G�6Ȋ���Y�X��TP��{7��?�KE��t�)׽�N3����`�swc�=�ō|ZT� �&�0E�bp��q��-�w�� �<�K�٥�PH��>���i�)g����}I�Q����󒴥$��M�RV�֤�8@W�h�6/:�9���+��'��1�~DKz�0�t��}�kr��|s�_Lr�=�=�ժ��eE2�1� ��!�L�jg�9ً����'�k�/�z꙯���`�\��Q��Z��8SWj���4����ܼ~����Lj�ɅhE8A��KYF�&mX�^�L�Lu�-�3�*  w�4n�\���h�<���Z�B��M��>���fY��f��&2��A�ak0MH�E k��B@�4e�#��kl�<E�o�ѐ�
��7Ӳ۸��cM)���F�6��f9Ϸ��%����R�`��- 4��2w#[��T���C�����������v�R%���=��1����x��ꍤU��A�nW����O�?x,U���Z4�BVy�f��~�Ӂŕep�!6�N�V�G���Њ%�\Q�.���/��,dˮ��|���s}��5_o����s���L�﯅A��ApV � �B��H���$-EJ��}���g\��c�����4�'{[��_��g�w�;��z������tv����n��қ��\��M-��S�f�2���wsg��x�i_[�뇞s_�;�����}��+'�������^W܃P�>T�)ȓ1Ȟu���[��G����N�4���#��Ⱦ� f��!nZ�~[�o�����x;�j�� l�I#	��FH�FI&�r�^�w򓍵:~�!��J�h~ݡ���L��e<��/W)�~�����<#[�_1���u�2��ۥ�݅�םJGE��l���EO�V٫�^7��A�绍̾Q����Mn�RLΟ� Ncj�%Q������������ M��o�� ���i^^Z�(س�6Lq���bˮ��=b�p� 籯(����<zi.;Lyć]5h��g��u���Uh�rK0���*;��?��y�埝0���g~�w���˰�ҵ��պ���\�=+��C�wg���$��m�幓���������i�;������ʻ7��׮���o�7�V�N�� E�MC�4�1��ps&�F�ٟ� H5�w�I��ѹii��� A�nhW#���A?��֟�:�A$�)�qӔ�,c���Pd�@�S=|��Z����R�D�/���$�Hp*F$ސK$c(�В�1�ɐ%�:i!$_�.�o� ��Ix�"�T�T8��U�W �3++�g 35F�(��ǧZ�i�p��	d\
��\J8�:Tcq~q�-�K`W�0%�YVdZ�<JnJ�Jtbz�Ć�@�F�T�G�������lF����f�]\�j��o9�{�-�w����:5W��k�:����D�WqJ�s	gA��I[��Ѕ6Sw���c���z��/�cw�R?��,,ז��Lǜ��q��t�����NhҞ�>E�u	�ą�xTI�x}���Y�`��'Ξ�A~�����'�G�>F+�v̈́������On���׮=�u��Z�A�F"ސs]a��4c�_T%9E�	�,d�����?�u��u�a[�\���	Or����X1�V��UG���eHItB7��nj'�7&e$3�\�H��g���}��\H4��3�d������͏@o~�MX*��(u���?G)ɣTs1o;�\t�zm>/ypۿ�GAi�,��|X�,�W�J�y��A�|�1����9�jVn
cR���Y��Mh���m"��e�V-"wˍ3׃�)�WA����`8�����Z���ݫ���yX�h�\�:ɲY�5D�RY�����PC����"�D�L[��P��,�@��������7��O������7��z��:#�q�P��Br�Z����_v�A�U@���4��p�j�Q�v���g�Wo|{ac���~���29���+[�>;0�ot~���.\���d�V�<����(�!�`�P�M��G�c\i��@&� �����Unv2kLp�F���C�����@ۅ]��������@�t%^?�*�3�m���������ۇ Ѡ�>#��u��j� �+ȠI�X�̂�2�.�6�"�"��%H�¢�E�k���4c�j�LX�L9*������������.s�w.y�����S6�'-]҇�NR��@6&�[�XX�k�=X;�75�]���T@E`�a0�u��CqG����g��VWW���<?��3a�� �a -�O��������܉�mQ�����-0�+�1�a �aP�Pw2u�3�U8;�
c:�	�Ş*���x�u��HKZYqw�|��W�_��o����O?s��5[7�p;��7����X����:I�YS�7[�A���˧�Z�f���ۻ�&��/�7�/�����Z�'=�c��ĕ�?_	����_�������7��F��~�-�EA���J�:���&��mJ�
a�C�̜�!�:d�2T?s�o?�a����!t&c��9�>2b��0�%#��a��f�F�N��HL@���{�I�W0L�/m ��!Rld�&���)yNa�FKdi7#E*X�ә��lf�Y�<0����l��$!��	T���:;"2eS�ݺ���f��w����&r8J"��ǥ�&Ռ3��.4 ��0��P��#���`
Z�A���&D!7�3UѸ����h..q���D2|���u��M�X�L�g�+��	{��)gahfVÀO�b"u$�6�I��<@��y�+��:|?R:E�&��O�۬c��G\kg�vo���w�տ��O~�G/ʿ��3�=dW���
ȶ�Q 2��.J�)n���n�7:۩���to�;@��jN��Z*5�N�7z�s������jcc��ݿ��U���V�$�lW�_�ʿ�}֪��ի�7����ܽ�����sv��*~���,���{����F7z����Q#UM�6��e�s����d:�J������� �:8�}|�	2�Ĳ�B,��0�fS�1��>6yВ�"5��j[Bd���&l�_���� ��Ŭ,3A$���g���ɂ��#޹s�gb�,��|��a,1��$11en�RKҼHK�daF�.��f�'�-�b�2f�m��B�ґr�0�wai��ـI"�>d�̾��2S��'#wIJ��"���s�~�E\�]i����ߓ����"��%|�v��AT!Ny7)ǷiຟVS�X87�ĵjM����вT�,F��g)�ǵ�����t��>u���k��'��O������'�6�ʷ�e�ޓ�l>��n,T��%-�\MA�:�$�Y�5$G�H�VA
`��$������8�JC5�*n�Kӭk���>�_l�j4Z?���я~ԭ��C��'4v����ڵ�֍��w��;���f����T/<���i�3����?`�U"n�cI��Vt��)��e)4����Lo���Y�ԥ:}�[�l�\�B�bd��Rd5�NhܧKАAT�Na���k
�^:�^��2�.#� ֛Ȝ�Y�6ٯ�O�W�.&,��Z�,��!��
�V�R�� *��9X�3\/K
��
�-�A4E	��C���w mi�.�rI��t��oSd�:�'R|�p��)�㌃�ߟ�a|M�������6� ��4�������h�*�U�� 
XV�aYG㙸S��`D)\�d|�\V�f5��-�&r�~V9C���2U6��47[|�w>�`K'� |;��21��f*j΂*�L�xm�:�W�2NUQ���2j������i��^Sot�ο����������=�����[�ه#�|�g/KY�v��`�H9�$2���s��+��p8QL���;�֜�rpppJ�>���+�j���Zk�l�.�0���wk�M�Z���c��V��+T�>�����/}�?���Gg��{�����I�N&%I�7v������<��a�w�f{dCcD�բln:����+ӂ�M�u
>���� �o݀���.��Aw@b~&�eUf�ĂdІf `j��ԍj�8�!1ꐛ-���ux)�_$�*6=�ȒI:��0 fY^T=sa�V��
�[���E���H�@������rՌ�@Xp�|K)}.�2[��B5� �YA9/���9�����RJ:/ ��d��&n�>&���^�
��M���U~�N��+��Ï
�K̶(XU�st0���O������߃V�ί���AU!)�tP��Ud����X��`^Htk�R�x��(Y}G������L5ϏDq S�f�)Q�\q��=,��w������u=�cXx�<D��s�S���״'�A��U�#�X�;�ۖ����`@�L�c�=^���"�y��U5S�����?ӻS�����l��G������ 1^��oBok /�T⦜p(�͋Rb*9�  SZ�6!8`у����/�ﵑ������t<�u������k���[��[�W�O>�۞��,�q��7-�jp�eݼ����kOF���r����'-����NH5=<sd��A�?�=AB���=��F�^M��Ty�aDuZ��^���Z}q���_�WG�p�~������ �:�/�أ�WG0��aGUg S_o��ƏlVF��X AV3� Vj0F��O뒢�Pb���
��#��R�Hb���)�o�٘J��3R~wI0R�qV㽋��m@G���,=/��Us%1V��ꔺZ�O7ƀ7�j���{%��?���Νf�������4O���s��������	����P׭�o�|�(dE$	!�#+��M &�,�{HPes
Yd����]T�� �b�8� )O}x���8��w�:�a�`��
w�$J!թ�:��,[�h�ׇ�677����+�ׯ��ko^2~��~�'�ϯL����ɓ���04t�6OB� JF�6p������dd=�J5�Rَ
$� �\ՒɎg&Q����ig�)��]��^�_�>��V�����ry��w�U���xu
g�x�'d�o�eL�~%��Y�����7��v�4S����Σ�aﴙg5E��,�Py�WJ���"5�(ݚ&�[(4V�߽ č�S��5�}6@��t�$T�Z�M:�Z{B��a��Ѓ�w`o8�A �'2ML�b�'�d���"�Me�F�AB�j!�B�נ�<�[��&��v,��h�ރޮ\��{�,S��n�e�0ˣf)��F�d���E{�����2O,��'!�]��K�GN]�1���tL��R�6�}�8ń�#+��G�����A ����Y��]����㣖x�秦'��a�̿j������=��@��1�vf";R�\���T̯c�����5/������j0��H����+koܴ���`#����g��H\��p����f��1,�m�);jz���w�Ad� b۶� �0)U��&�!d."3K��?���o${� �\�X���XF�z�������������pb�A�����r@:�p/<�
��Ѱ2�vQ���ƛ/|�=���H&�R�ygS��M�Ī�K��,b�B���i@ݖ��U��͝$�\M�f ͩ�M�Vg�BJAJ�BȰC�v�j{	��<���ן��:���_�W/�.�c��H��2���������ƒ���(g`A����K�z���نD_ċ���5d3J�d��ø�x�����e��(:i�S��|��aH��G��$��J)2~��t�C��0X�`�U�m�n'5�=��8L���M��'�{���I���ǰ�{t���Z-�]f���pF�18�*7,�&]�*G�w�����ۯ,�����5-�ǧ12�a$��i�q����h^��3��.����@����c��/��B��n��o����?s��ߟ�������8gOn�+o]���<ϟ}�m+��v��*�ܱ�cN�q�-.#�hB�9��i��"c���1Db��XM���F7��f4bp�Fn�����t�֕m{g�y��c:�vs����|eZo7�f�	@�k�������1[�ꆀj"���,������}�>��S?�JY�9�ys=�W}o��$�.KS�=#}�\��# �H^aQv���R�\�dEd<T�Me�lb��bN�������f��զ�&O�yk�����ӅW~������;��xڂ$|�RgBTː=ժoTV��c���Ԃ��F�������!UC�
L2��lc$]b�wR#�s�O���9���(�G�ݷ�_�U�:ōYR	���(�$9><V��j��d#f�T�� ��.�-d�.~�r��bV�Z���,����cmdwx>�����C�lu�8t��ndQwR�9d��P"����̕�ʙ"􎩑�d�����>�M�ߦ��4KT���b}�`�~X�@�1Xd�����p�'���������9��[��ua�ۃ��gNm��MX[X ���A�?�TQ*!���2��,���,� �T�S�H�$����Н�Ȋ�����W��dMBЕ|?��t���ׯ8�9�eedW��j_R���������U���Ս�ȍ�;���%���R��R�����̣5g� ��e�����v�0T�0ԇ_�j5������2~_���?�Z�x���i+������,�c[�d�B� '�p$�[x��FN�;6�\bSG��Oe���+�ҼA�C��8I�@UF�a����Qm�3�Z[����[7�&���y�Ex���Q-�<���������l��D��2f�8�Z�@&+ېj-P���TV��6� �L��.+Y���*��ҵ�	��������+K�ͧo������<;�R�1�����$�T��Z35�B�`�������X�����T��� ��_���
�9�t:N!`���nA�VA����]�;�S[t|�sb !9���V�+	7[q*ˑ�~Re�WR�@a�8b��A �;]g�pGnST�&O���$<�Q����͖�h?&� ۋ������_�(���.->��;;Ɨ��}�F֟;w���gasi��W`���Rg'I���69���n�4�K��J,����$Q"�C���I��K(¤�"I�Q]1�����B�!k0�̓8��C&�L��U�����q|���{�n�>5M{��+J�z�������/��e��KMtE�r�4�<��#ix,�J$9��HJ���)�"!B��gIb(y�_�٩h7oV����{��(��$�d0�$�[��Y,*YfhH��<��8�ZQ�ؐYJ�@��q�YP���5��w-�}1�Cu(<�Tw���hx��*;��������I+�07��z�zݮ5v�v�����=�Tk�����߀����/_����2���S��p��Uk6�U� +��D�����M*������ћuЪK�d�!�8�DV��O�=T'Kc���ȕV�.��{��1}�5��9���1�ϕ�Wl)�(���QW4	w��'FI`K�:��iyn��๊�#���ȫ�,�h,kg�_%��CL�z�!<rb�-dm�{�R]|����+��61غt�H4փ0eCI(1�&�A�uS����٣�y�)��;D�᫽q����B~������[3�M��e0�l$��O��a��h��m�_?qj��_�����o�7T�3N�y)�=��_{.�����5x#�Ϝ>	V.F,܄���R�w��F��)͜"�x������&n���\*�ș��̋yD�s1:W��_��F�U�	JvK���A���(Ɇyg��)#�$���`�l9RݗE�	3p��S�1����3���O����ʤz�S��Y�I���,O,9�t�4=K[��
>�"F���yfP_(���&J� '���`������(֠�͌y���W{ ��a�ld��dlM*?$<�'䆎,�"6�O�]��k�<:�����曋k'��p�������YZjN%�;O����o�~���k."VAu��2�񄔎�CX]_a�0v��+)E���+1Y/��:T6 ��۵@����*��9��4��թhZ��xxO��`�_�]�ǅb�w0�1�"f�@ l�խ������:T��0� �� WM��&��W�>�;{p8��O}
�=�q�b0t���8X��j��s���]P%1zC*_��|i"�$�c�*T�l��e_��t��X��,����H̀
��qo �εYZ�������r�9�T��up ��7��pc�1�~�V�^�y�W��6V��׿�_�����(F�-w�C�-;7w�G�]���mx�G��'7�E�q�q}ؾv��k��~� k�Uf�ԼAݗ	�I�
+��	6�c��hF��}�v��n�HF��"�N\ꨔ�4s��t�J4�!�lYXf�
®�麙'����O�2��Ej��"d�z�$ix�i���#�L��{��H9	&Qo�*�FVj��5��S2O=)�yE:��5��|P*j���>��&���$P���d��YȰ,6��&�q8��¢���\XQG�a�%�����=���{��D5�����������ݗ~�����_�^�����s�T@ft��|�þ8���aG�W6n��*hf��B�H!�5v�!�	����R�n�jB�����/ҩ�.Hq�ϏY�@c��r}RAƗ�wa�&�S�в4-R�G5�y5�y9ƲI�u��~��P�F��A�9q��Nq�y�������tLq^�&�NX�	�G����Xj>;:�._B
����M���|- �=��Y����I`����,����аH�8��Q�2���b��w�k�.tY0>����>t�kT(n�,�t�A��^��E5b�"p]]Y�`�c?^:N�MVАц\�M�gQ�f�`�U���<��p��h?���zp��5ߐ��K?|��K����f��)M����-/�y�*\t]x�?�o��5x��Yx��)8��K�&�]�<\�x(n�8�:I4�6�*4x7���4⍗jI�K5/��+����Ki3��#��4��M��(b�ҩ�8�F�F���'r��W��B|n�C����}���G~~�
;Bԑ�J�g��D��J�H���$p-A����M�68�ѐ��:�Cf�0&�'V��q7\:u�Sܔ�l�\7��X���;� �Y>��OO�.�rb��[յ���8��w ��;�����ſ��7���ϟ*��h���H�Ǣ��q����?G���b�l��B`ULd�)=�lV1��5Ng�"D	�;���If w�S��@��p4��t.>�ʯ��,�3n�!0�}�+��s��k")�TU�1]_�ȥ��ܔk%�����(e���o�bKr���Ѭg�&�K1Td�������ZDpu��V��l���������ex����#3-�-�;�Tx�,���{�R�����{Sh���� S�<p	<��5�fG���]tn)آy�r��S��vef{H
_�$�)���P���ي���c����B�i�W^q���o�|��_~qD_l��?��Ak4BF�U!U{���.����u��g���Z#y�PMj��3�LX�1uc�)�WELI�p�k)�Н��C��W���("�m��a-M�m$�������A|�%R˿�C�KQ>���!��{V�}F��pKCP��(�n*)m�|s!�:�U*!�Z�Y)���'���]�/�9~��u�+�>F���.+nĐ��"�ߥݝDsjC�^ S�v�S�U�?��>���+-.CD��v��V�����+�n�������۷�������C�i$�8�Nx�ִ�?�q��"�T�E���Mv���y1���[�\�`U�D�V��A�X�dBY���V��n	��F!��o�`��4�@Be������AfƢ����]w�b������/1��=���/�M�����S9Oo�]�2�S��<�Aa���84&��PcFt�
t�0�a��)<�n�z>L�.�ϛ+�.����둆�e�ch�G�So�����{����~zp&Z���g�<^�������mY�7$q��8b��4��}����.n$��1��~p�����(�ړ���%��E��7'#n qps������'�M�jÙ�%8�nA��6�n͊�adb�x��ㄞ����Q�Ϛ)ʚI"�WQ��(�2w�JE�L0cEH��$�L!�bY0�8M��j���S��D`��(>%�/�5�8�g�o�	x�l6���V0*�:�1�ge�XY���U�U1�=��H�L������ԩ,��y~9����k/��8u�^9A��������97�T������W��{/����'A����*�����"����T��������P�e�	s-��O�4"��d|�|Y��������P���ᦖ���1�2��3����1X��H^�g�A*4�)5�I��{��c����5��ΌL��[��i��X+)�����e@��e�i�Z~K0@eJ�R@i�&�ƚ��� �`��S��n��@غ�v�����	?b�E�YA��	�a�8y�2
P+�\�j�" �@�Zl,.��X�^��t��0�c����o���{���� :à�ܒ���EG�R|n�
�{M��rC��k�_�*T��z������{߼���������~rIV5I�-duV���Ȟ.u�ЙN���>�1�"��Xo��EXDFA��$�]��ɘU�b��#�����@JiV��Pʍj��^>���,&뷒^/���B�Oф�.?K�:K�T�&��L�4G?��͸(�&������ܕ˴�$/�7����dnj��k©U5�%u�A$�Aq$�?���mO��¶j�i�K[��O�47;ժ�t3g����V�e��җ�x镟o~���g =�ɉz���"���Z++<�C�.t�u��MڝL@��1p�!`��@��Y�/�H�Bg�M%4�j{j���hWA����1��н&]�Hg"E�O�.�2%�W�=Ii�G̝��h�QO�̳Д��T�Z*�^���|���қ���ִl��w{���~�U�:_)U���cg�A�D���~:���'��ެK��:��{����VU jE�*J�z4�{^����<̑~���ќ3Os4�nQIQ,�],վ`_r��=|1�{��yxDf	�R~��yxx�{�gw���0M�򕫰��1�M�0Mau}v��蝶t��_\�����3��S�Q������ٔI!���./FĜ��5�T/,�Sј�|�5����p8$�ok��(Rt�p^�uy�u\�+c?�����B���_������v�ޣ�}8 wKx�Z:���u��7�/B�aJ+l�G��8���.N�6ltZp}��O�9�����5p�Ǖz����T	�	E�N�'��I���(?�����D"@N��f|�hѻ��3�p��C?dmV�\)�+���m��Q(y5R�aW@�6� Pa�\mC�5��F9o�p�IjC�VΤ���7׋mϝ�g�{���7���ݠ<X�5v;�.��k[��qfݍ�)��^_M���(�Z�}q����_��k���_��W_}��Y�^�̒ͰV넜��( N 0�I\��Cn�'�p .��իW�����ڔe�'F)�S���=��Xa��!h����ǜ���"2W�9��+�H�pq�W�C�)e�f�$J|�S �E��C_	H��?EF���B���h��zdl�*���zR�rVbOs���q��4�k�VyD��l��si�:\8f�GMU��t�`��j��1��ُ6�-�;�s���������4���(�{�,�Ů��x�
�^����	��q�׽:���w,[Z���Ӊ�KUV���^-�iYT9soww����������?���M�����ƕ�F�5�L�Nr�T8��w@��q2��Ng�=܁�E\ͯℱ�`�ڨ�%ޕz\��ĭ  �IDAT\��B�7������p�\+�l]����D"}�	�Tt��QA�O4l��o՚0@�;�<X<S95ʏ��L}�����t�y�ˢ1ڊ<�YS�b�M�È�~f�cj�E0�Nmk�S�T�^ߩO����s��뵙S�uq밻�1l��I�_��V�m����Jmn��w��Ӈu��g?���ǟ�уޙL����/&Iܭ5k�u<V��\i�P�X#h��,'���V�=�G8S�3Ug8���!I"9���=�йp�kB�]��pҍ��d��I��pQ#,MTo��q����Er!�ڍ"~7�`,  ��wY���N��bL���(�a<R-1�d�|�-���sʪ�B��=)����_��@��C͵8�I�w��YQ��PkvXU�������M�x���!�*jk��x^�Y.�k� ���"&�e�� ��Vm��
Gքk^߰�1N5Q����sddRνw��2)�n� I�Q��V�*���:^�0���?����~�ɿ}����ͷ�����d�q!��ζ��9�S��p]�����=��La2M᳽`!�8�l��@�����I��lt��F��澹��6��Џ&օ+T�L�C}��|��8��	 �=M-!z�#�]��C��J���3:���v����!���<ǗDV������t�}�^���ZP�����w�?nw�wl�y�z?\]Mڵ��j�'�	y��w�f�<�<�?��w�ٸ��~�o��O��a��y�΃��x�i�[kA�s�k$y�6p�@�d���<!{�s�E�,�we��mc�NŶmUl�v�۶m�b��vr��]����}�'��v�}����
k��I��^�
�s
\V����*���1;�����Ԛ<kE0r��l�!k"��IUI�b�^Q[^
��T;�\ �lv�𼈆��U��7'��
�P��-X=�n��?�}��ج �B�]+��ly>�6�e���XSb�f���~q�Q �	sʸ&�t�C�+1���HF
��h�+vb�|�G�Or�E'B���r���x�i8CvD�|O��vk�J��@ػa��j<��7���H�`R��t��p�~�1���ĽY�?[��X�76>�z��E�]�
e���A�r���L"�����[��Yc$P0����f.���:��Z������M��Ag��;lbG F���\1"y�:婪�xD�m����Q=����h�O�s)�`��K� Uؑ��
��V��3!`G*�L�Cb�c>Ҩu����-�X��~R�Ǉ+��?��ȉ.�_o��e�3��pخ��ki�������Ð@53���ٻR��	o�d.JϟB�Ԉ����=O�u����rb��c�%Aّ�%���� 5c4PD,�vda�.A<�Va�?՛�9�- ����@��^}�_O<�%9L��� ��i�ʵ��ȭ%"!5��*Ҏa�^t�e�	D�I��e`t�^N�Gʀ#4xF�z��r�@i�������aV���T��ⶩp��v~���d�+��|��YCH$b>I�ܧo�����LU���z�k9.CL�N�Gl��Q���}M����.ٻq�]4=!vc�=G�����d��f��+!�)k5 �-*z(E�G��Fe�.,V!������k��8�'I���9�'\>¹ ���ͻ�B��).7V�Fq[ɫ�'W� �sw�`�Ĥy5�Tۦ��z�P	׿�C�Y��tu�sZ�� ��6���y�X-�U�!��sL��(�����x��o]���Y�L��Ĝ��Ȋ��M�.�ɕ@қ�^To�h*Nx)�� ���wh�wh'h@wS"9�BL�g7u�g��,���ٯ��>��������%���/�_@���Ϸ��������%�=�@�I�i�v�"<*8V�hCUY4CA\6:�<�v�r��H:%�]RR��7G�@ɝ$IAS�!�����y�O��y&U�EI_�W ���1&	=�~b���j�{��˫sU�k8'0��D٬���/�׿�sܞ�Sʲs1�v@�qGz��k��K��f�
<��r���ֈ�G
����m����y���^�������z;\8]�2ę�4�+�\��t$q�������Z�>R��u-"~S�+1g�>|��Lk�/��a�b�0�'����
\�d6��dqT������=u�oo]�	1�I�F����?9�0sE���ҭ�-�βϽO"JZ�A�Pa��hKYα��f��Xm)d���;A\��F��v\q+d>}s��	��
���E�����V��������m�;6�)W5b�a���c7^'Ҡ�kI�t-ع9�3��paI���ۺP����b���]sm\��,tZ�̝�r[KT1�P�Q��Z$���b{��O'Y�䘐-c�L��!���ņ��u��\���Q����M�hy%:�1���P����Ӗ�w�����ʎ�Wj�����2O��V����׷�����2�V�/V�_�P�Ce��ù���۹DQ�+@l��l�@��!IV��2�D(��('+��<Wj:��r2U�_K�U����ӫp��ET����r�^��u+��<���u�n�@
��<Z��z�_��k�&�?�*�'�l��*A
�M}m�ޏ�=��$G]]��9����Z�����{�H�7�ck���&���҈g�����Oj�1�n� �N�O�<Cƺ�x���x�����1��8 l�N��[ń/�bG)'�"����}���"�����a81�C�M�^��Z����p��	�޽�U��M�{&�^�*1��Q�y�����B]�6�����!��a[��١�)Q��3ծ5^��Z��{m�_ާ>��蒔]%Vr`�-�^:5D���ߝ�>��vؘ4����
�B*�o���F\��d��y��M��L�Ǯ����b�]�x�}|̨.n�~��{^�l�M����)'�U��{�� }��	D�Gt8s{S��9h����}w���������.'(�������h�%w�#�{0)�	H���/)�x"ї��� ��X�6eE�H"��Q[�)�	��e���ϻs�_Ze[�uƋ���qT��#��#����^裬va���:��p4~X&���
��[�	ߩ�nCn9~4��:���	%:ݬS���rk�P��wo<���=����e�1b(�Th?���]}�U0��pj���ķ5'�[���	Kk��X����)�����'z�үʝ-������~Wˋ�v�w���Qy4n�
�J��(�-4�l��ft�`�9���W�U����^-a%�����ZK1t�;��B&[��^]��C&�[#�r�"9�㳨a(
��=�7sdzvt���O]6WH�)^F�#e��/��.��,Ŏj����Z��ԍ��wc�d���4�6Y��T�?�¶O���!`+��!�!�n�PЯ���?n�K�L�
����!�5ݗ��uj�_�C�+��>�~�g
�\>��\�D�]�w`��#(y�i����kaɔ6���'\F�ǖ�/>�]���Si��ӟj��(��ȧM����5��W�@@�Ka��<����4�(���
���Y)�߽_�mؾN��ѭ*J/G�p��p32�0�^1�1�=�YP�h�:%iTP{QFJ�[9	���S��Ж��~UeA�F5��
X���E�U�Lt�.�{�U���K�^�֧��]�F�~/��ү�H�� И�����3g?)��7>g��>^��ڡJ��f�%q[�ق�f'�`���
T}V��k�x��)R���-�$c�B-3�3o��_�@���m4�!�|�E�N��=L��c7��Y!6ͅ�Y+>\���X��|O��J�On���e��.|���^`�\��L���H����4�����2&��}[u�WcN�\��]@��fY�{����7 `~��`c���t�N�c�Ki��o���|.yM@o}��6��?���|��WF
d�*|��ρ}���������ݲ�������l%t�/(5�h=�*%�/��k��f���6����s�ͨ��{�70���c�.�<^�	q�@�j����e���z��K���|�,?nP��m1|��i6c(#�sOJ��TA��_+���2>�zoyhs��>���K��[��$J�6����כ��"/��߷��/��<�׽��`��rN�����㿼����я��
&_�w�ι�(M�
���8�h,�ݛ��w]~2rL��1̝Yޤ��!�g~̄�閜�B)��P@���!�>�'�k�$c��.\�َU�jiNUX8���F�dw�}�@��Ş�dt�����8C�?3K	�I��E�6������2�s����d��p�V�[�/B�ԪB8�z�5���'�EH�9�况4'ne�ʧj���*��V�`t[l��7gry� ��p�������f��G#��ws�I������V�t��0�<d���u"5y����b_ X�(�����,"��������s���B�!�%Q�@}��GnQB4��Go�oZ�� �Zɕ��,�(�O�OFw�&��d����qy�U4��[t���<�s�V֠�cF��Ɇ���^��)�P��?���¥�<�|��/�|�	�{|��y$}��E����}�ۣGx�*m<�A�[u������Q8	��`0��izmuE�+�c>�A'�(C�T@�:F�އ��А>�Z���X���ɒ��#ط��r��$2B6;zV+�W�F�6ׅ��-��~�O=J�rrFMx���?�KTiV|$���^o��	gG�
�v�;nw�Rw����-���İ��'f����a�M�fu
���~�	��h�g����u$~��]��{ְ�##�w�t[:��Nq�V����(K��Y�����n���Ia�bh�}���˒��Gݜp�yW�*�0�"�m�b�Hx��H�i�����	F�AͶ�J�R�T�VI6p��j�d��
�6��C������M�N(jzÉ��ë<j8�@]Al�(=6��3q�o�kZ�Œy�[���b�	�
}����ڱ�����/����s&�:�|���T���9qZ-,1F=ؒ�'E�t�T�r`d8�]�r!/�F���
j�~�9K�*��f�����@_0����ɃWN�.�Y�}p�W|�'�b<��=*���C��_&`��Fb,H&����{;�Az�L���P�^�����N�~v"/]'��R��Հ����W�k]�=�In$�{!Ѝ�j��:U�$:�b7����^���G�J�d>��g�(LY�~7AK�u�t�Ų;/D���=�A-�~t0{����7w6��{�I<��[��y]��!K_����/}�Pfr$��2P<
�L�G�s�5�*w)� ��M`΄� �M��N��ȧ%HnHC�������%F��8�H�b��ǣU�xy����g�J�]�֭����?U=v��9.�/�o�%\�bg���ҡ��X�Ϩ�Q6r���-���Y�S�t���~5��ٰ��+���ꬸ��fY��� ������Y��o���P���c��v��3sD����Bc��R1�R����y�J�fZ�!#(�5��k$4��AC�iac��U�ե�;-OgrzUt�l�������6�`�$ƒ����LG�]���Eҫ���
{��%�(��\��&ֹCߧ�	r�҉����~�X�,�И�q��i:���A�Ľ�� 4�[k�#?�Eo$���s�1��Z�����X�Q��e��_���m`����P]d����z�Kn��PnO_Ucnp���cE��d��1m�kw�.����+������V�i�c�V�k��s�K,�L�h�gG?���|�~�-�#�yϿ=-@~__����0l���G���>��.��p+��?j_�	K2q(u	�|�Zf#�.��e�
`!<I�2��	�C�M�t�\��ՀV!�8�E��)52k�����S�7����z�r�s.-�Bsr�,
�4�6a�cT�;�s(h#�̀a���Ύߓ�ν�-�<��?�<���n�y����r�i��U�i��sR��5ok�FC��r�\��D�����m���vKl�҅={��ّߨ9�׭��s�ZB�P�\���i��,E��c�s�(u1-qyΐ�>���3k|�eC��!�A�NJ���J�d5�Bͼi��rVQ%J)��л�B����`<�����A���4�}ǎM�G_���غ�/���z�͇��Ǐ�b���^����S"�GП�"_gFP-�D#��>{��40��ԁ���r�����~Wa�(�uS)�yy;��ʳ'ؖ�{:웧��J�h��AŠ����pܰ��nNlZ_`}��@�,��&����� �}蠹R�-�[� -���A�J�m������5cY*G �NJ�8�C+r�7O.O��r��hp��U#���ӯVYk�?U��ð�qN�����@nwc=�(\q�����o����$���r��D�m3^uk���\�g�qP.�e;漻�B�	TS�����RN�XB�QD�d`�ݨ��z�F5*W�Zç��z]���i5�9�]-U�On�e�E�wdM*�� +"�:�Y�Xϐڏ�H�3xJ��=4�׮�+��~T�%�,{�'x�5��� ����Ž=J6C�t�4^p�&�V`����E���|���Ɲ�ܛ�e��	{^�I`�X�J����	U�c����4� ���KB�tƓi5�g>mT��*��p�>��/��מ�l����k���vʳh���������f�
u���t�)0�Ώ���4�s	;]ws�Bi&�\S��΅	�]��Q�|k�Z��o�k=�vRh4x���qeATQf��	�^S�1UF��ۢ>97V�: k���NM�W���;�yp�C��3��G�E��C8;6SGs����u�j�Q�������ش����,>TY�J��G,���a�Ҳ�x�]K�P������l�G�"��wn�>�a����DP��:j�8��m�f8�Si$�l�2��0b�:�s�.�6���R���#�摝.��ft�ku�/�~j���_����8�ș��G������{7ݧ]>����?\��#���!�P>�����u}-���l�9E�W��!~��]�Fd�x��͹�t�֜X���^��s���g�����6p��j���Z��gNJ��E��Y�W-�:x|��xn����k�$h���JR�Ԝ�����èx��h\��zS].\�pm���54U���$��C�+�ȧ�ғ�D9�V�a��&:�2<)t�gA�m�3�$�fnҥ9t�,�"(p�2��&�=�G��(,��t���i�Z�*uV>}� i��'��Z�/3��J�`K�O�� ��Ӄv��=�N"�T�ZMȜ)V��]"�M]o@m����-��>�����;=�o����Tߣ�����2�C)�J?���	h��C�2�z�	�_���e������Xt���t�۰��|�}�3M����y��JŔ;��JS�P��&!w����Ӝ�D���jT�#�Ѵƪ�5@���UF����I�ܹ�Y&h��?�>���2����;��m=�
���T�p���\Ѯ�)�L�JT�N�c��V����{��ƾ�PP[Dy�n�x�;k�4iP���k&R�+��D��\M�?m��?楽Y�P|�{q�&L�y�����E�6md��+���/=y�K�G��#Ŵ�Uݟ~K��b������W��V-�����"M3�������*���T�L|m5?Sg�c��q2�c�]=�����B�;5���8�ް³�'�x/o�inM�	��{�a6�dm<�]�L�J?�8�.�$�]�Z �	ٯ̍4��WR$�tƟ��\}>�!��u���������a�S�
Vb29��!3��ad���`�F�7�:��I���x; I��Q�	�S��!y�_N�r�� I�y�4VEɣj��?)]�u����T%�(��щ��J�l���
��:�.�Fw5�H�4}�@sKHZ�S4���E��m��eL�!2SЊ�ȶ�sk]J�9�ѝ+��岔ޗ]��e�����콙��`v�ȇ`c��ۯO�:�\&n T�E�Qǧ���~�"�������� �"���p[Ӳ���z���]s[�o������V�	�9��d���'�6K��3s��p=�x��R4�0^�u�2.G����%��o�j*~Ht
�ɶ�y��cF-gs�Q�����	
 �c�Ho�VP�LxtGW(o������n@�����ԇ��f��Uٳn��~��pʬ��9�H�\��ZFWrcZ�"��s��Q�Q���9����BY�I����&gx�0b����0��-_��G�YY��ڃ�e�ѫK���V��jN���,S���h�Z��֭Q�o� \rM��0*��u��p,A_�o%��OX���K�i,��	�-�hji��U���@�|=��qx�Ј�9�H�G�_�껠?�BIz�e`z��h����;-ʧ�Mpd��jr�{�tta�B���|�ޑ^R��܌���N�Ǜ/���41��|xk�&��U��oy�OUڽ�1�y޾"5�����ދ�+$遑��	�����!�j@ϩ7��j*"��纽����R��N�׍&�8-��R�R������<KPHw�{P��u�k~�<���}g�DF�sb��!B��HS,�M����T���°N��k�Y+VO�� ذ���l���by#�U���$-'{מ��-Peؕ*��XŲ���$�)tq�q�V���E�zu�,x9(�M(�P赙??��t?Di�r*��0�-�����7�^�r�Y8V��KL�0+��L��ߚ�D)Ư,o�(�6�CQ��%[��X�{��@�6x+����d1���3�z�տo/� ؓ�� ���f�ףG��9BarT��@���8�>T�a[\��Uf�7Ve-G0� V� `�����5ݽ�>�HT��	�J@}͈QIZ����>`U�T<��6{"��3kV-c|*:qq`�B�]�]	V�ه_�QSf9(悔���v�Y��RvѤC�{���9.�Ϛ�x��SNs�1�I��M�3�o2͏Q8Y����ū� c�h�̔E3W<x6hR�ܩ��S?�A�0'j]�A1k��C˵ED��n��퐡��_?Y��&�F�0����3��*Ľh�D��+�eu�c$![�e�K��<���(��7z���HY����",�l-+��&�jh;�wO�K��j�ӛc��|���]���M�������PKq�iE���Vu�c
r(�E����3�T��Z�$�I��"�C�wI��~i��r�KNp��5�~�1G�RW�/V�a` �"Y&	)r�|d�;BB�[�H/Y����"����[M�M��V�}�c��fh�߄���CW��d���wO���lrт�"��]v�E�O.j��X��W?g��'u@����o;��bM��+�;ra͑�,�K��)��;��-�u<��CH1��	�X���:n��n�v�;�J�l4=��኶_ ��ғB\~L�49 |����u��1�A�sc/�!���~����[���{�Z���x���_�rZ�pe�3�k�l�r����N.��-q��Hހ��W[y�c� eftm�LO��$o���ez~0�E����Qf<�L5ɫ���)\B���	�.�P߿��[0����D����,�H �7 �]MAx�G(Bm��[r�u�
��m�Ȃ�+(l|��	����UT�`��4�_�����~_�w�8ۧĔ��d�"����@+B�	��"@p#�Q�_xV�jP�(.�MȽ�J;3��K�em�!�i]���>��ZwI#��2�2�z!�*��p����Ë�ݡ?Mhɦ0��H�x�GL���&�v�n����!''����*8z��Lj	��O*�/�\�m��a����c�L�|q�G��N:wjĆ_��l��`�OjC�%,�	'�0�5b��������37���5��9W�o:�G�p���U?����Y���ؽ@a,��J�
���1B���b�|>a /H�G�Q���6��o�9�,���z�MQ�Ŷ��O5�5%�Ņݽ5�B���/u�e�՜��
�}�UJ������K�Izg� q@	��ص_p��೽�v���:Xv����'x��Kd�V�9�*��`�Y�A	�F�]r+�T�Ƚ䟬��=d��z2М{�K /��Ө2�q"��TG���i8̑kqf:5���qt^�������>��Z8���ZW�� �R�7|"~�E:bm��)������D��P櫭{�|�ʝ�;�{���nFC�uRq��A�}4)f,׈wb��hy�1)�3r�*��?V�͋2�8��LLa?��~�6��O����ę3���L����XLuR�*9��r��w�"��kp�9��Ä��KJE�vP��w��\�-2i�ZX��Rm.�<�Fs�T��M6CO�a����O�ѳ��ik��nIf�|ʙ��	�&C�g?t�[_z��?�Ъ�C�#.	�x�8����f���fL	Qk�{���AXy��ݮ�OPM���Y���`2�O{m���ґ� �=֎,�|�4��a+��~WMʭ�T�r��)Z.��~�����ŤWx%�QH�ݦ�*��b�q�	�� |�h
��-�W�B��3�y�7<,OC�5�?�`+��t*��GN_Ņa���{`9��ڋ��%$�#9 ̩���ʊ�^Q��С������nK���@$x��"��3�'ou,�7�ld_��>��Yv$��_��ڌy�z A<T:��c�p��i�-١��/<~�{(�>�Y�N�AT5��/ʴ��*��@�}CC��������7����`_�%���PEP����1���v�J&��m
�CBw�c������T� =��Ro�a�4�Ŗ$'��K2�@I��,�q �[p|U��p,�H.�Rt�����{�Z��F?ӣٺۙ���������t��W�蔛��c�PPp^�@�7�[�>�,U��G\�_�������IX@�K�6᳊�Y���~R'�cҿfS"�C�ܢB4��V\Q��������a��U��p*����R�P�Lf�-��A&Ѕ�^��ʳg�I��*�ω�"�����Y�a�q��&r:3i�i��m~s�G޽��̊���9v��/�����%���"T�4m�>�mQ����絴6������@P���-9�h����#��T����%�c��dʩ��p�� "��'��+�L�R����:aQ��$��I�4jk=0hsf	 q=���ʸN�k�mZ]9��� �!oް�^b�Y̪RmD��b�7z�}X�apj��sޤ���_� &r�i|�vo�0������K*��)�z{�K�I���28ta˩y�̧���ߗ�������ސU�vY���M�]��6�ch{@OZY3����Z� !q�����pH�u�8Fz��<,!��i ����2�0˰��lx�R-U���8��� ���h�?{r4IV
�J����+5<����hBL��i˅����i�Y�6�Y�
��N\k!�JU��@y{/���26��Ez�o�2�/�#�TK	7�����b�6��U?�S㧁ja�Eq�!qsO��S3U&M�mt��A�xG{9�Y�����>I�2t˰ah5/]��׃0R����.4;3�Wl-��(Y�R���Q6�.�l�D��ͪ@��[���e�۾{�5���T���N[�S@��\�`����rU�3��r`�e���Z�����I&���z}2�K9s�U�v+��c��V�b7���r�9���ut��=g1R1>UE�|V�"�8��k����@������x!|$�4jh��k��ۭ�����Bb橴�צ�R�k ���EBI	;�;*Z6����=|\�Ϙ��:x�=to�%<̪,D�+q%��ܤ��\�А~�������g�����bW��z9���AN�R��yX��Q�~ˢ;l�(���h��uiz�z*ɟ=�����mj�3Y<���`x<�)�$u#��|3�x�/��ݬ�QN�ҡe���h�Q�̢DR4(h���,�����P��		�k���.
Xq�B�i^�g��-��|���[VHH���t��TnNz̲6����t�g�,~0�H����}MV�x%㸤������㎊����AK�'աj��U�"@��#vg�M@��q�tE�r�~�[��y���mvBWЅ*t�dX(K1¤�+kL�/��4�Q=!��F����袑�)+�x�b.�?��p"�r:�YvJ��Iw4��Р���I)��
V~����'��ҁ��K�B�^�e��s�+/%�C�l�������W����*;�O��"���Q���q��@���0�f0`v/�p5�r�%��w\S?������y�itg��?��"
)4i�g�Ԩ����?Y� i#�
�p_����1����X����j��osi�6+�
(pc�lH˼Kq�32��i��K�� k��y�0R�]V35�MO̎�!���	��&�[!2~�[��!<�N��_���R�$jW����ŝ	A1��dޒ�6�f�>�++$�_��Jν��ڎ�V�V�#l�D�6� ��o��=��"��5i�]�DӼ���l�>�f92~��^ͷ�)����~1u����:��}Vz8HC���^�� � b��y�W�;<�9�e�u&>�Z�Z�E�ο��&���;]���u�����c�
G}�"��'L��D@�����!�:�r��/;�5p�	V�/��!�
N닟q8��ISYz����(t�ngޖgO�P�S����k�-~��|.���H���`# yZ�j���	��x4"��D����{o�z��z 68�t*�m;ש�|�=�?���98���2h2���!R�π�M�=�?��\�yL�$�8sCu� Za�$��4�MJ��L6b�̒<�&2��j�����^R�C����X��+�<pNטUM��^B+���	��v��,��GG��҇OU���=�l�w�6��(K¬�C�'�� �p�I~3c�e�
1�p(�s̻���,9Ml�%ι�M�夑3�b'�J)7_X���"ɔHgR��8�RJŒ����Dbr��C��~���@�֮��
���y���}�������Ot�g6ր$������� ��t�i����j�yl��$�wP�(�ПO�Z֋qh`U�wE�ц-�i�	�ed��o{6H��,T���j>����@�V֡Mg��!dۜj�)���XU�Q�0*D��s|v���'���A�Y��`��mi�6L5��Y�p[i-�FA�6��� /?��-������Q�d
��K��K��l�̻ �� af���gdSsĳ�߼��Ec�{j&���q����~C�L*]� ⑧�F��G-zm0GF��u<�+0�=Ἦa�$�i|�(�P�wRM�K��O�@Q&����8h�2�6m�r�35�g�<�N��v:�P���[��_�4��F�ڵ��5 ����-D��v˝`��]{���hhJssƚ<�S)>�7�o�����!����
j>�&Z���ւK�Q�9�9��V�)��Ĩ�֕���1K�۬���n �0ț��͈��@lw�a�TV
#$$ܶ�8{� ,m6�2�K��NL���@�;-xB�dh���3��)
P��<Z',��ۇ��1�3mE^��kNF?�}
�?Y
��#�85��,�;����e]:���"!�s�0��f~�l���O����\�����x&���������X���0A"	Sx������M�dY>\��.��!_u\��_��҃,q\��
���X��$�'�U�9#$���9�|��
�So��^�|=BǦq�B�?w8�o�i+����)��E@؏���^�������|��R ܴ)!���������%}Ȇ=�D�qڼ���Q��@ٙ�Ӎ?p����M��\2�~mS���'��,K!�d.��o-�P$�D���RP5 ��ى܋�F'�
�O"��&�ѱ?�＄�C����\q� ш�ة�[s�&%��m��t��4���W�ShT!�8@?}k��b�H��+�Y韃#��շ`�^H���A�({!��\`�;}츄X]�sy��i8)���(I�t��?�(Ko�jb}t|�!��{~��/}�bFqi���f*H!7S��A�m9o䞅3[L��7o;�@)U�8�{c�7T�a�W�g6i�G%�@o�)2�2�Q3�-�V��-bf�\WK��`���;�f���L�U����
�@j��RN�9�4�"BmNm�eJO�k�dhAmI�s�@�/	�DN3<
b����O�A�[1Vp�'�[�o*DK���fm�[�n
�+g�0�^/�� �u�p墣�ĖH���b�U$�A0h��j��W�lJl'~��.�����j�7��Xu�
��3ʽs�����耻iF�t%��y^�f3#����%θ6�M�%/K�,q��On�U��JՎ{T%$�M��f�*g�^e�c�_�E���(�S���r�4~�k|M�����������m���kC�/܈���Z��X��S��.F�H�:�>.�c�k.��˛i�EE������]�46G2�fKE��}љ�[6y0+�LJd��潅���+�o<D7�q�VE?��$�7� ќ��7�t�W�N�]��9Ŕ#�Z���I˝��	B� �/g�:����q>RW�^�j!��f`��u���sC�h��b�܀s=���	I�#��^�.?R���L��c�����7׿s��v+BjW�G+m9p;���N;�=X8,�|���NslOuϵ��_=1�%��x64�+ć/��ɞ)�<P%z|x
��<�q�#vRY2�	��Wwo�}����Ia����ב��O�f�N-mOV%;-�NjFb�1j!d�¡B�+v���X\�G��9
�_R+�$!/��U�u���(7�K"� }}�+E�X�����b�_]_��������_��r��@��XB���1R��uQ0�"aw6`;gP��g� �qs4U�Sp���M<g�#���=�0JZ�`D��A�����r�S��3q����	��u�(�uz�3! ���4YG����n:���UmI۟�Q��s(�Lu���5#��T��]ʏƆ+�]��I�����}}����Q�?ܡ�㵣�k�]��2�������������(19P��4`2c���n"je������}k�*-��͞�M_����`�h�%Q�~��2K��6H���RV0�.��O�}q_���|�,85��$_<kʯ����s�D������%F��/o	Tml�>�b�հ��w�u-�l؊�R��ɴ�'��*mqz��:�R����7->��b�%����������z��LE.�����������
@q�ٿ���(��s!��eA-)��)�����b���.����ߐ[|Yz���ڲ=�	$�χ]M�m!oy����V��pӽ�Pj����]1Y�^9�9a�ej�`O�D������
5�:��'%^���m����,e_49uZ�7��,�hn�$�<2�$D��)3j���hk�%�U�w7���'��
��/�4���=B>䮣�ܦ�Q�.�dK$�K�Ƶ8%���w͈�׻���I\���ǒG���#-"= ��lix�"/i��T�e�&*C��hG�tP'o�8p��V�;��Լ"s�@��1�h��^O�|?$9{ �9�
�)�<����_�l�K������U/�%�_���pI큓��z�n�r�P�rʎ�������
�1���i��J��ǐ�[����6/qA@8�c�.c/�K�����Y�r җ��m �- ���c=���~ͤ�J�v�]}�� ��E	�m�W��������{G��A���*����9C�q�Rȟm	��!5���4�@�tܓ߅�IT�k���n��|Xf'6+��QY~C���!5��69�������:0wA�|�'y�L,�G����*D�������0�m2�5'�rfp��P>_�0���%���xEV��B.(�L�xı�9��t�iZ�s�TwOHϹ�����Y�Scw^�ښҙ�,�&�]���M��]-�Q�!*�H=�%��H�����5n�"�[9R徹<�;��������U���T-I��erS��	M停Ql"9*^��|�A���T\>��tީ�u�g蟆B(�O�9�ݱw�_�n�Dp HlQ����OO&����'y�Yy����N@9s�fi�R�+J��uQKx�?�J�T�`|fS>��O�n$�U�v�c��Lӟ!Q�ĭ��.��C�^_|i��=�<�ጠ��V�E-
)ܭ6�o�N$����lZ�9&���u��u֥qL�32ٿ֎L�����j���E/}�ݎ��_z�\�$�5L|����ҵ@F��
�D���%����_.���Ri@��hZ5Q��W�FeP�&�o@0T�T�(geW�\��:پ��	D����G!�L��W��[�.-2��	I�٫
�M�=Zi���I�x�N6�ζ�/[�֨�,��f&�P%��0�>k�T�[U��{dFy-�3�9�� k��(�1kKȱ��@0�N�,�y��H����|�6T׊>��E�9�Tm��o���a�A��Rꥰ��!{���P��YD�$x�19���&i+Q�J�K�������@QQ����a8���|T*��2���|r����M'���tS�C$�ڸ�Kh��;)���D�ʛKr�|	���:�A������uFy-�D�%�<o�CϦ��},���~�,�䫰���bXa=&͖A���j��]��F�1p�G�䧎L��M4B�J)<��sC��@���xR=������2�����9p׵�]8�m5�m�Vc��mc��Nc��v�vҸA����������5�a 7��~��֤2��W��M|\gAh�����6LH�R�~`�%���.�.xa#���\-9Б	�=�P��P�=>~,<��}�:aA�?(�	�}�[puK��sr����Y���?,�=<g-.�è���ЛQ��XԴZ�7��R�菋6��7���A�R"iBDp95w�->�ꚤ�]�׌;���d~�#b8�QIe��<�Cc *DT$I��ɱh� ��>n�f��3Вb!>$�_�plw':Z� ���I�q8jO��Jh��-�F޼���2��C#�`�%��gϥ�Y�a�{�-����gx�o��{����[��1�j-�MI�<���	ej����vLs�.�H�{W���X/�n'<���7�z�,CeTJ��Y����S�i�־wD��J�gtDb��3�4��{T���p͙��O	e�����3�cEn�5$�����.�fd�g^�P�Ɍ�걇Eފ3 �lE��~keBk�谞��J��yce̹s�W
(KC�PL���D ����k��"	|���߉��l3y8�Z�[;�U��DT��'��,�:2�o�dx���[�f
�#����/� �,/Sݡ�-�9 |&��[+E.�ԡ��ς_N�D�%d��	sJ���p�K�4��Ⱥ������ڳ[�˓�԰��y�CRѠ?M��1���h����
P�7�7n�t��\��j/OJ��������p��AN|����J��!�5\ѓT��7ŷ�VTܽQ{-ܷ�9t+oΌ#�Et#�t�.�������F���N�芘q��Z0v2b%3A�3;&w��5�#G>c��M��"pڊ\�.�'a�O�����@��ݧ���݁\w�|i���I���6*� ��L	U�|�7�sUf�MM��kt�CYd��]ɬ5MB�S�ti����($2:�����G|���粘 ׃ۜ{�9�7�������BY�]w5��ВW7y��G��ɗq�f�u�ѢV뷇��KC�æ���B�PI2��n� Ț������G} !/R�`�l�4�_�;}� '�7��S���c�ΖvzN����&�I:;�j�^|l�f�\T�ENi��޷ВƇ$��/G��9��a.�4?���E��o��:��n�vdĬ��GN��dG�b�s��s��Y����fp:5�=�x�j�S��7x6a\���l-9p9b�P��ØJZ��lEv6QXan0�R��Ƨ��Q�4vb�6mx�%�2�g��IZ�ۺ��*\����P�4k�L-H�VD��X��m3��o��G�c#ʚ���U���:3�z0]�U%�`�� |���\\�3���l絤�v�R�2ت����¬����a���H`��E�?��\�ZцN��y���3�h�N�=_4��V0�h�H8p�m��8��kq������'�"�����$l��/;2$�,Es�G�:�>��~����ӫ8���l��i�ay���,)����� ;x��#�V�{z�`��|n [??�M�實��5���d6ܴ��* ���(��q������>�j"GaVV���Z�]�_�h+Ʈ\�K:�����}g���TM�@���������b�ny�K_��p&�rr���;E%�I��ѷs$;�*��[��eW�VJT��r*��4֥��b����*IRL�-�&yT�kN�0�{g�gh��""\��v<~�M܀�_�� V�XOZz�[�؁�����\�m���� �/���C���ۭ�0�G����*�N�(�%��dYT1����{������)�%{ᚚ�A� ҕ�h'c��-����̙fÕ<̾���%:_��BO��jh�5���֔���h����u��k�U��-��k}Ogн���q�%Ss��_i���'�ni�Q�N� t�Ty�5���M���ԉr�"O��ij����D7� ���l
+3'�k���ӹ;	���I�5(ns���PW� ^
�M'�`[�A�Q���ē<��9!a�IEB������I������à�"��Z)qX���ZL�]Cq>�&n�k�;�����W�}�^��n�<:��E�Y� �ń���>F���K*����o�8�E��K=m����ƹ=�^�����qq���Rh���?n)��x`:�9�����5_���+��
S`�{ɍ�m�ڢ���5����Q˦���m�[f��T4?�*���I��0�S�5sf'U?��h�:�5θ!�|�Ŗ#���H����`].W�ֶ���ɜ��X�¹C+wmL�?[���������Ç&E�p���I�����M`��	,$�:�l�\u��hl�Ģ�v��0	v���Xx,p��X�0y�M+���PL�k9*b)4pI,-:tso3bw4�G�X 9Z;7]��3Fb��fo'�)��<Rl��e�hܢ;���������M����cGqL���ȳ�:&��xJOK��`XH�Q�M��;Xۺ;�*�c02�w�	�G+��Y��#�&h��=d�.������]	�>�"��_�z~y��]�w����n�e���m7=�<|�gړRL��}xz�/t��,<Īz4W���v��G�t�.2���uPE'Z�ZE�v��rԿ������m��暚!��5���j�~uU����}b�E���+`eL;k@�Um���\^li��5.�5i_1�����;<i�%	�j�e��LB����ަ����2����Lxg�w��EjXw"������і��PiX	F�����~����;@e�;<?sB����Z����(�O�oH�nJ��6Ԝ�h�=�e>���h]��ҥvۜ����n����G��hn�_��`�e|\�{lѤ �Ô(UE����q�o���/��Y�&�u7��j�����g=L���1b����L�� �Sw���&��z0�HŚ-�Gu�Ƒ&`��zڼgo��w�=�w�]��!�A qԁlZ"RA�`�:T��XǰK���O^b1� L��] F3OP��6��OFCT�腅�['+W�ǌ�?�~ާX����$Y�L���к����W�j���' ���.qOH�ll�#H�yǳB�o#rʌ��p]us	ć3 �H-�JG�6\+l�&�+~��
p��Gk|S�$tQ��:�����ٿý���F��<�8!��Β�z�a'������š�7��pB��>��)��;�,�CÃ���(�^>�u��<Q����Nq�"Fm����ܰ�� {�P`��%�S���Q)��:g��}�i���!*>S���dG��#�����L�1�6O�.n�)��Ŀ���V �
_�!��ɼ�����M����2H���䧘�U-3�e�ٓ��7�Lp�>"g��lpj����W��4�q���5�$0�OzUV�
m�g�LƝ3�n��©C���`��;�m�j�+�t�L�7߂7@m��i��h& 0f��p=�F�`�%2�)��SJ���Of��ܠ�e'D�Z����^�=�������d4���p/("a����Y#`٨LP{*"!r�sU��6�.���ê��I�q!�a|W���.^�_t�g=��9����cݿ�]�G�ɷ��Pgٕ�|��Q(��.�5�;}��Z%��لݜ+{t�/� �
X-�t#8N��]^&I��6�=���j3x�Z�� 9j��(��KT��ޏ������"a%l�7 8���Y�h�z��&AMf�Hh5O������?�,Ec��hs�<_\ሄZ.5�X�o����2݁r�ӻ��'�	�V]$����A&��C��L�_��{��%sdY�in�Ȏ�9�X)�UA� �����k�m����
�t��`�����Ϭ�&2���\��/<�c�Z(�cV�ͺ'�/�g�/X�{;���\y�D��s�G~���,s��J�����`�Pg�Xr\	BX�
Q&��^A�Y=ʇr�����_�D��&�_KD��&��e�7�Ys8�ae�&�U����f��ک~q��A�n�+����Wz���V�0�E�h�z����=oL��@��Ԓ/�F!/0_J�ݻ��f��KH�?S�]�d?�i�E8,�Z��mIs�Z��_���U㤵�Wl"�)v��ټGe�S3x�ON������Vn��u�ҵ�c �N��YW��!#����pqu�I�Df�۲�p��G/�X&���(\��Ww�����U�~rZ 8T��`�� 0ۻ{w,���'�a�;�hA�j�����Y�J�^�&���� ����~E�D��A*E�kO6�_-X�1cށ�HjQ�)��N>!).�n�Y���5�NV�{�u��B��B�N�%���e}*���Hc�鯊wZ�d�3:肠*�*�����2MZ�����y�΢|���g��V��ɫR#n�Z��)�0�ag9�$X-��"$Sn9|�g�9c��6��{���M$8��H�hk=���|��'��wP�sP�m��v�� ظH��'�,4�Z�)2��-�g���%�$(�^>����VX��(������O�؞X�v������-כ��f̮�瓗���J6�xX�#F�0\�y��v�N�a?\XHմ��7o-G�sD9��~K~���
�f��$��:W��Q��7rn7�g�o:41Y0I��jn�Òݸ��KO����\HL`Sk:	���F������������̒t�b����d7�d�mK2�;P���3��V�����7�/����xxlCO���*�uɬ�Ab��n'�������Xw!*z����H*�	l�^�*A@d�b��\�`Q����f(Y�Z��a��Q�[�M�8��e��p>����6\��ׂ�s�x�T��}*\�bᑛ�}��&n���w4�M>���[u��D�P��H_���yZkJ�X��X6�!�/w��5���j�6�h3d
�� �㼁cmݐ��7�CM��,��%n����!kj��|K�=k�Y���1��sN�N���`(�!�������Y���Ҍ�]J��B��s^�����4�tZ�-��-�4b!ҺQ=�h�/(K���mQ����T5��X�!��'3W�h��)�T�k�����,T����0�q�b2P3��(�џ���y~�#U=[���15� ��~��� 
���t��q&t Ax����B���҂�4{�vjF)�{q
����H�r���	MXq�6�Y(�ی�#������G/�BΓ�s�Ï��²��o�3��O�\�?�JF�)�~�&"Ξ�MbɞF�f���.	I\"��du��[)��ͼ+��%X?6=>�XSS��׷�����%1(��v+�%���P��Pji�~9�G�U@��-y�k�Ʉg^��W��P�d~�Բ�����=��l/6٦�B�D��"��#ܑd+
�F_�*W�-��q	Y\>/���E��#gt6��.n>V��+���O ��r~�đp_�࠽hʕ������I`�+B���6�+�dx��B�{�[DE�@��E[d����7k�G��5��"Fg�Y��u���x;G��ٝR�	�zx�/鶛`V(b/ػ���� h7%�t�kXIe�%Ly�_�Y��+�g������r[�HfH�T�A��=�
��3��H�ƖЍ��g_��Ô�%Z!.�SI�\�fz�*�f
P��NmߌǅxuÅ.AJ5��%)ϧ_ǸGcqHA����wZF�#K�?ҷ�[Q�D⃋c��+,R"�?��ePO�A�~wg��,Ȱ/$�i��V",V�[>�B�D��#��R�Y�'.g����&Q����1)���-WLʛ��]�DuAe���q������),�,�Gl��j[@��pΝ9��Mp�9��c�Ҽq q�2(�,tY����6 �Y6��6rFҋC��'7T��_���>���𯲍z�J�H��4��T���ȁ�aP�~i;h
dP�����sԮoi�<�?a�����N�y�VA�Ť�����8n��I�^R�ub���n�9f"��T�u�M�mx��B߮�`��"q$��?e�leyº5�?�L\`T�e�Q;a�&���pKO�h�)?�/��O��N��� h��9�Υ��ԙ-i�6���="��R�b��5A�^/�7�+���%b�	���o���a����Н���w�WQ0J)t��C{�_ݓ�{8����}E1:�/�bH�zW*uAh�"|����C4rr�r|J5y��o�k)3��n�7��ҽ:��'���h͂t]���YO������y��3|?���h�J����M%I���"2����%�Z
-�٥#��-|+����b���8�(%NJ/�ys;��	K2{�iP�>凉�3cǟ\D����>;Um���3�%c��{��OW��hZolx�@	2�>����ݘ>J�
���$�~#t>W��c��\���:]�4�V��� ��F˵�#���0��r��iJ�X�?uۢ�m���ӓq*�X�0-]ն:K�h��B*܈�V~h}�b���gwqsH�����QJ�y�fU���ζ��@����1��λ�3J�5��
�s�t��~�s�\س4�o7��W�L��]�]��ə!��Ó��Ӕ���A�YS*�.0�$����Ag�&�� )����n�w���5!x����s�D���)ځ=�j{P7����A;�dj� �.P��j���~�_v�U;5<:�����xƣrAI%�����~&O*MED�$zuK�[(Ҕ���6�5�<z�#?��0+S��������Mc{��!��H�"�p��$@��v{D�pb.��T���ہs-�R����'�6����P�Yy��}{3?T�(q�!���N+�
u�L3�0GO���+ޓB����:((i���g�S���}�KblΆj,�L��$񎺆��6ړcy`|)��95���w #�7��Qz��A�W�7^�@���m}Ow���3&�L��|�ڊ��]
X��V�
~V�Y�#!��m��{ҍ&�X�ɯ�Ϗ�=��^�{f���Z��=E��]5jF��i�1��r�$��_����M�ҙ������a�&���ӎ�z^�7���sM���x�t�pu�,��{I];I����^r}ڡ�#�
��\��V�8m���d/�4̼i�+DonZ������f)�=F��޲8�JܼEd^�J*�E*���H�,�ˊ�M���^r� �����~ɝ;`���&�����>54E��xظ�9G#d�������&����!�=�L5|K�k�H��$�?Z�^#·ݵ���d ����J+��?�ň�O˲�ԙ>S��`!ٸY�!hN�t,�(ΜL���s2h|����7���!�c��1���-���q8z����y�pۧDE��_�J�Z{�e,#RRK��QN��	���^�Cn�(Zzu�S,Ks��<Y�i,����bMs���Q���=�MUŧ#�N/� �n��.���g�b�!�]N�JQ��+���`�E ��&C�Q�{+��#���S/�GI������#�U��%H� �0��է�;��PFo�:oB�c�cs����Rz塺��!�t�Q��sJ�ۘ�q"���p�]|�`v��2�"���p�N�Ps;$��\T�Rմ���'d�Cva܉�*�֌bE����3����Tm�o��׈�%tՁ�<��嶳B\ ���e���˥-B��-m�b!�;�(�e��^]a��A��F��A��l؛�����c������3N!"4�}����&�_?��^���6�h
�H�oȢ[��^��Qq�y��M�q����Y�ٳ��������j,�~8����plJݗ��\3s|	Å�ƕ�k�Om��9NN2�V�]x!�6�R q�]��5�1�Y.�%���9J�&tƱI5�SY;t�I�P�[O��팅�0��D�\Q_�R���9ޞ���U�Sj�z�=��@�� .�P��>1o��{�	�~���O�b*5�@~�nq�K��=l�m���'��������o��]RZ���5�Ɲ�_�=u�П<~ oe�v?�����A/INM;A�Y��T�6��&}�S����f�F�����&���T>��Q�����?��Wz��$	�\��j̍��_���׀��h�����x}E�y79�ݘ��QO��
�ͅ~;&�-�T�KA3�j{�`H�j8
X������;�.m:��yJ��15�༸͕oLz�re�j��{k��ه�dI��!G����)�P(R0=��y�3�|1^d�F��(��W���_����F��!�[�ݖ���,�6�p����qHVv�׶��4�G��b3��E���83��Rӥ�Th����C!{n��J*-��-�����S����&�ȩP\�2�>��4�h�m�������w�iI�T�"����M�{�3¬Ψ� �|�����Yڀ�j�S_�����#M�������\���j��\A u��+#�)���qJ�{c��[Vn�������\�x��Sd������v���2�A�;F5�Ӆ/��$��ԁQ�"������%����(���ot��~ov@�](��`��?ػ�S��f/X����TV&�����u�aʤ�fb��1�cɬ�kS	Tq�,bH�:�Uq���6Z����u��sE�ڜ�9�Kƨ���4e��z�#�����󀩐�2��A���g�3��6�K��o7�t����	<u$d��KJ��Ԃ'��.j+78��^�Ɠ���o��=��n�ʡ18L.H��vև�ϯ�v\��{�4��n	~kj9��ʋj��������uh���\>и�O�ݙ���'	!���%Pm�ʰ	���|���<��ǄR����v��#P�qk���N�I�B20q��w����{�g<�'׃�b�2��OU�^��Ԝy��sl��<���e�T�_�N��������Q޲f����D+5���T�����3�)���_ɑ���-.)��N�+s ��]�4&�ɬ}�/���y��6����:� ۺB��*N�bC#c���NXW�Hy��Q��*i|�$*�#�<8q�N�P���6���v��"�!�vb�MS�#6�&pJ���L'ٞ�aE;j�q�|����kXh�m�nQZ$V�Ձ��N躝�cʜj�����c�0L�ֶc��t��ł���2Do!�eR�4�H���b��X�u
0��[�i��d4�Ύ���ϙƅN�_�j�@�(�E̲ �ٓTjyz��c4��[m�~�tP�����ߊIQ�~���Ye��H`ϗ��Kdp���"?��t�\����B*����Ksy�1z�:D�?:���{š����^@�
xe�y���=�;�9��|�<�IL�V0 p����f��	��wb7HC`6�ב�Z^�1mi��s=����r?�tKn�d���M����z�0��1k���]��4�n�\˨��������H	ӥ��6�
���eـ(�/�g���z�AI�tt��h1Z��j
��u�ĞoL
���?7\eOt�����:�?��'bx�"G'@{4*��*,��Xx@j0�}��d����w�Z�bM�v;��{ɿx�������W��2�����nY�e]f�Yt�6�"����(�t��C��x��-� ;$����h���*��Ā+K�o�3c���iCG24�vU�� w�Ύo���Sɂ����rᕂ8�?���$�V~�a	�eĵ�Y�d>��Qw׌�R�A_�Nzڢ�k�QA�z����P�G�-b>�Z�#�r��҈��1�M�z3����ϼ[�^��̙z%���@Ls��gUQr�s���<�Q��Ս�3ܒ�bLAo.��t�Zc���o`�4 �0����E̚�6Z�Y���&@y�q�lT���@0�~n�:ʹ��WԩJ��!�J��*X�p���z<�5�5w��n���G�UIL��mo'�1>����m�}�wzdr|z22��i<�s��őn��r����%�����t�oa�tf��8��	��"��Pj�c�	 �Ӣ/W	�Q0��A�ڽGnz���:?��M�iSW�=[ȋ���L���w�5,�0�g���Ш�j�~[Le��~i'Sow�8�� j.0&47쁺�b:N&���dמ�ZZ�Qs�F���p~;]�5�#�y�V�LaC�md<�"x�$eΆ��ث�f����*�D~Ky�$?�Zp����߻#��ɱ'�n��`Bp�&݄��)̺��-�.+�JC��_��f�0<�3}p���Q��3�f�S���cc�Ք~	�	]�̘4����,�w3�ߧ����B��I�hȸ�Ҋe�S:���:���j�������%y�Zގ����:t���+�ł�0�qd<��mJ�t:Ғ5r�8�(c�1����A�A�U��!}xT���]O8ru�%anj{�i�.i�'T�Ta+�s5B�=��$aF�̆�[�t�IуP�kK��ٹ���(�謨��J��]@�9�2���ms�/7D�>��U���)���� S$��T�5�=V�����T%9�t�h�}X��.�{J:�ȶ���6�RXC�}퐬��U�]a%BAN�����`�!��,ˑ$%��V�A�)��u��,�J_ҵ��ՙoR���-�3���-.�i.��Ic���f�-��-���^Z��e��$��:�(�Ol�
9(4�
8o���(C���{+e���r�����k}ט�jU���'hr&��=�kF�S�m�w|�6�2b٥�[?a�Nıt�8b�� mw���5~Y{:��$bG�Fe���*m�Þ�x�
5:8�8�F����[��\�0F~sd��'�&(y��av^$v9[��V����o��
�(�֦���8��Z��IV!�N+�);3L>����"�:#݊<�5嶌&��$oz���O_���x������O��$�r���A�y��QДز� ��'�Z�@�n�<�����?o���i1{f T9��n�Ew�/���K��{����eaP�a3W�d�ʂ֯�`bpz�:���,�QGB��6��B*�b�꟞�
8Yd^fǉ�M�<��ؙ������r훓�BBq���Ӻ�gũ��=)j��d���B�W�H��g����?!iF��|�:���	��t*i7����6Zд��y
��̓�nl���Gi@���8_N@�nDo���kc�Q�
3ɭs��n��	�ћL˽��RQ(�>ɬyKk؀�7�Q�4����/G�;.�BŊf��o�.jm����.�x�㕢��t1�do��B1��X�׃lt�Q(�2{qo>܅D���MNf4����C�ܥ�6����b'��	�>X[�^���
gg���~<�b�U<&f41/�b�V�=�J��?wf�a�������;�%3�|�)&�[�u]oɖ�Ԩ���Y���/�(��Z�*M[�/�|I�T'�7 ��1fscj������Q��&�����c���6���V�N�4Ĝސ,�����X����Jݵ��p���.KWb�*�!BfB�����w6}��D���5	:vv�xD�8B���8DjF���Q�a.���38Ut"��Ƞ.�=�O��*[')^	,��u!`3��U�w��d3�����òz;��Uܖ]��-X?V�l2�f�#b�.�:�퍠c�i!C��Mo3���(-�@���qRvY��#��#.��(G@�����*l�bV�]/�ބ���va����QLm9Uu\���4��!���D�xÒ
�RTi\�ϙ�D�G��=Y��i �Q�㚶��H�%��U�����ɡ��+�4^��4�dv���_����B��V1�񆏜��R^K�[D�g�Ū�kL{

sK
��Z���2�"��|m��g��0Њ�&���A��w�X�6?o^���Nү�zm:�RuV+����-���
p\���9*���TDz�}��\Y��#�
��|,�7̼g�Ы 3�[��n��~��H!ޙ�[�d3j&zB)ƅ_r�Yq��]%�l��G��G��$�#ej�}l�z12-6)̗��k�!kIܱ��X
����^�8 T&��y�
Iy9�j�=XEyk��'m<����T��҅�0t����m�k�m}nR	�Q�1	���5��d���K��n��l�#�8�|K�����.$���[ez߫�ג7�Dq���F�^b��D�b�r��X�����mS0P:S�*��ڜ��e5}ֈ�F�� Jel=n~�ŗ����O�L�m�6'�hXQ�6/���_b��?&�"g������jp�o�"�
��i�	ݚ��5/Q��Q̅
�*�%^�޾�VG]Bi����^�F��6�# =�[;��9F��m���f^D�&�^����DS��uX��xlƻ��ڶ�0����ޙ�uk�*������QbZ����!��;�/�����u�1�g�@�s�rk��ρ_�c�9/�m���]Jػ"���|%�,9������뗿V�.?�}'p.�u�.��2�&�c�␷��.��
׌Qg[a\ �:���]p���x��������G���3�/V��{09	/�����6�t�5ZޮC�Mg7��"7��!g�(]C�A��$���rOiӣ�Plf�t����D�g�� t����N��-�	��lʔ��x��CTg�e�"���G��&�W?-�~�Q^&6l�8�w���^3�oRJpA�)z�烎F�HY����Y����.��c��)Dp��om`N�@c�VZެE��-Xb7����`d'Õ5��
��r`�9:2��_ko_j�����^��h3��aw��Z��<�3�i䨜('(�%Q��r�0��yG�FyL���� 7W����߯�T�
h�YF�4�r�A`����y]�����i�T��x�b�����#���j��+(�~j[xzuR���Kzj�DM��vc���r�h[3)!�ϡ��l��[��_���@nOtXE.�%ߐ�^�����}�)\���ѯ��rrxd�;~Xۡ��f\��%l����M�z}��d��0��B�U*�v?�pZ�O�r}6�諸���JE1�\U#��!��Vi�*�@H��7����I��Oy"�Z�gYWf��Y�tX�	��j�n�]�!���4~բ{�v�}�1��^t���X��t�Ѱ�dX�W�u�nUf���H摾ا9}`g�v ���X2��:lɤ]KЍ�¦��T�W�4ߡ�U�:�n���۹[�pY �\�p�3�u��%n+Ljx�]�G�����f)�Bi$�7��9����[z���V<��xq_�EgL�Ε>���T�M ҋk�g]&�#-Ԁ���_��pXG�A���2٣)����n�s�?�BoM�-7��-���-��6B[��f�9���S}.��z��֍�d�7�O�N���!	SP�sҘһ�c� �S�4QԿ�F���JO�p�AAVu6��F�ᘀ\ VD9��V�z ��32K4Ş8/� ��kR�S�B��콬��[���;�3����Lɮ��4@�96��ET��}*���<}mޘ�{P������E%��a�?Xd�Q��A��5ps���AaOR��������R�8��&��D&~�w���i4���o��Cg��v�@�}�hz}\T!���X`	"<hA�Y�w�W�Vŧ�B�_A9��ߝ��XX�{+w�bz��:�&�Ĝ鿌���2��Ϣ�'�!g
�.�#��qT�&\2��� ;���Q���ߞ�
�D�`�3ud�lF��,ڀ���L�6��f�-t� 
g ��q~���86^2ӷ7��C����מ<[F�����eԧ�1��^ѱ5����-N��(�R��U�_���H�����B��톽��Q���]|!v����Z�\���Mr�	@Dy������=�3��i����(.�8:����Zh5ϥq$����}�h����)����f�1��X�[�*;�����ڝj��1���5xy,���FB��[�+���Td]�T�{3;+&�)G!Ҷ񜮑����WQ���^�^����i�Rt5󄦐O��#E��6�^f�>1����U��?���~1|�%�ͳ�;ѐ�Zl�T���\��lHl�A?^:wOp�#u�,=n#&�����G���/�F>6 &
�]����L���VpB
"����K���(`L%F2 Ǘ�����:�B,P}���Lc��q�T�`z+ֈ�!kL�u�c������<����*#u��Հ��D�w?oԯ�¿�Fc\V�;4zs`�E��=Qg��}�98�����?�ب~����3�pTU�+����&t�{&��ǟ\Ŗ�	cReiև�b!��B�
M��0)Q���_
!#傃T�|�%#:�f_?"��<�c�1�����mԋ���j��X�����C~`�����s�F�����Z"6��I�X�IW#��P�D�"�~�nJ"�|n�v9�I�� �=�G�܍����"�<���=A���&���~��ui��<,�o�i�򞚮aG�H0��
�mXH�V�U{�-��q��&��5���qR�U�C&Mv�ҏ|V�_�M��.��NA��L��8}���ÁF�e�v�����5����.�R$DEkU����xu��"3�Ut�>�W����~�[���Vρ��hܗ;��ܧ~&�Cן��~�<#�ƙ��]�j����X<�NN�f�bùA"���M�z;�ဲ�٩7q� "
Dz!�F�3} g�暠��5�R��͒���,�l�Y�H��mŠ����|��pZ%�<ҟӒѢt3����$� ǼU2.�^����Y����p�<�x��Њ]�`��i���UY}��:������a͘'��-���"��y�T8[�s�C�	<�ѽk��'�����*!�҂��G����te����_��"�I`�����TĄ՞)Z./	��!^	���`"��n~<v��Ρ�.<<��ՙ˄[T�3%�C,���3j�Z g �����M��"<�Bk�Ϋ@�;���DP�X����؃9N'���Q0���a�-w���=����_.���[^��z�jP:�i�5ɯO8�z�/��żctm��k@ ���υ�r�o'Rrz[4?5h���nf�O?aQM���[YW���`�>m�V�lz�l6.�v���G�����}��E}��DH ����K��@��9�����&߱1~�w����J�5G�U�MbNg�#���I��
狞��ƃ����hm3O�J`D�v��N�ߌ5�[PЈU�օ�a.��G�R��9�V�")G��f�#�p&29�#ͬ�!�Nr�u;5�sʆ���w	o-K)77`��Bum;
֮�!Dm�B��qBˠ�\�u��\��D0j��k�������.�]�A����Qnb�n�"��!]���ś��G-�CL����ي�ۺ���߉?�M�&a����8��8�^�)�,�އ�ݨͨH���എȶ���`��q��şI�k�$�(��%{��~h�.��⻺C�����Y���i���Z���P��������A��U��>ee�I��~�Ղ�������(#)�o|e�H�.���B]����'�ȲQ��T7�	��@�x��튙,�.�%BM��F#k�K>� w�U	{�1�HO��r�`��8�v�N
��%�i+�}��z��a�.�ŀ���q���o[=̫	m3xL�&1<-kA�Q�C����=E��Aț��`��ۈrn ��lW�]iB����k����O>{p�m]&��P;��9ގ�_��6T�%t����	yKfz�8��t8�ʈ�������#M���|������a���Wvk��=~8�v,�FO�6���*G;�9y�ι:gG�u
wIDej�"�Ǭx>��ձ0�x�μ�Q�K¦�v�;�n�f=�zKY����?�ȟ�$S���'<7Qx)˚�2�:=�:%Ӛ��1�q��� ^����s���;�K�}����aA��~w�� Z-��C��է��>�e����	�3�̛�i�6�C�@�u>n�SZq���:w�g@�LZq�?���V�"�r���B�jD�����qajs*$0�$�E~��ΠF��0k�\��F��&�&O^�f	�$�M"���ӓ�e�DW����͂yެ�u�v�C�VL1=�Q��hT��%�2[�u|��*��c�J\��C�&���PZ�+􅍽0cM��B0f4�)v���/#{���>F�!�V�<�߳��~$ڋ�$:��՝aq��n#V�7�T��u��c�I*��6A�c��-{����t�Ҍ����hۮݨ��&�m۶�ضm4��d�Fc�v�c;�����g�ε��Zǹf�}1���D�A��*��x�:�2��4?'���ݟ>j��)Op��؊0�Rk5�ij�u�l�j��z¸���w��<_3��>m��:
��J��i~;[Ұ�EN���H�A��[.�'~�5~cr Pd�0>OW�X��<�h��$MnԓP��БAo�d�=�f��A)� ku�5�T��<����]� G�d��!DS�b(�V���Fq��p���k�u�\���S�r$&������Nn�4)�g��!�Z�v�F�gF���덏Q��
3Ӂ�AD0��},�w jW+t,TE!)h{0�6;�v�:�/��VI,��$(�W��`�<ͮ�Fx�%�d�kȃ#l���[��Ѯ���ّ/�e����iDK���l�P�&���xG(�{z�8|�ͽA�l�;QND��Q�Q f��>��ז{>������LO��74p�=���R~�Fw��O(g�v����Kz��J�&���ܑe�3�R��_HG��OkD���\�5�oEl������fL�;>h��!�Zv��_������A?E&�v�Ep�`y�[��*Or�7C���g{�sz�l��v����z���\��g*n:Cτ�)��qȐ�D"�3��Ͼ���@���� '��0�`FMU�G!�"�b��n�#I��0.1�8�1����I��I���⮤�Ӂ�5�F=!��MA����䣣{��Ƒq�&�oE2o:��M��,��� ��;v�0��_)�ȡְ��Y��
Q���$u_�,��]�p>��{:sA�qY9�`|���>��E�g0��k�ZP�U��o@.���{m�.׏������u雝�o�7/fCg�y'n�_tz��_�~߆KW̚I "D����g�h���\�2��>Oo=��_߾>�?Y߇j?p�V�X#��=��H��3��9?҉�;��Rk����*�x����Y��?7f��/<��K�4�y)���2�xr:��0�\�Sv;A}� 4A�=��I	���lAz־Ȁ@���Y�T�oZ�yK체fl���e\�P��(�5�y�Ïh{m�y-�*x�j�U�ǷB,N��%�jE������ ͖���I��t�'����-����L�~ZG�m�U���J�i�\��.4���7���o���y��%QK�����V
��ӿK�ŀ�u�Ґ�BG,X���2ߕ��#[��� ������t)USJ����,.�ym��G{n2`�p�-����)�&b)UQ�!������Yqx~+'���A��<`Ј(�AD��x� �C�V���e0v�l�A9<��͸�a�R��J�7�#W�`0��a\]���B{߾
�O�4� �R9��QQG�`�fu ��lO�'犤<�bjQ��'uP�ř~b���x�ka��e>���(��,�-�j�#��}�T6U!���I/g̺�D��un�h��t�u2\�\��g�7:�	x=�Jɇ�I�;)������?r��&:Ї��G4��čg��1QG��w���:]�LBں���H�%��Z��~\<J(�lNaK1��;��ʹ"F;z��Z��ը��K��)�f���9��C�}ŧj$�X����W�q�d��rX���;m"q�4�d��%�A����{u�z<Ю�.��?�z�0�J�D,�-!��/������ش�EI�3�ѡ�΂��Gk f�Y��G2��|[=��އ�!Cm��C���M��y�d7�I�4fP܁:�D7ú�z�$�Go� �v�M'��/��Y_铻GqڴC��X��g��0�F*c�������i��>��?��{�t��og���]4�P�&�g�x��-��@�)�.��iF��ʘ�$Sƺ�����U��_���3�����v!j�)��HL���d ����y�e��3Ot��*��x;�$�i��>/��D �=HBC7�Rt%iUF(;�P�[U�����X\���/t'�b�~nHV7ɪ�q�Q5���&� p�5ټV���8���m��>�Y��^��Ѯ�+@J\�=�R��8��gv&^|��d��D�4��)ܘ����� ���(�_@�*C`�p�_�������,t)���((���	|6�$F+�� 7��\u݂0���͊�e\�X�[֗]൨QVu)� _v�����Y$��ש�&ʂ�l�+�գ�F4�p��L�1~:F��'b}#߸f�\�L %�2F�Ku�SV#�����/���ik�ׁ.C}t;ėM��N� �1�,�D_�"n�c�z@
'"8�*sJ&Ԯ�`������뵀m��3�����Sn�=�:��k��ߔ^7~"u�T��e�X槊�m������O�	oQ�eݴE���Tԅ1�p��FG��<t�Q�nZ�����)�{��H�T�Z�X�S��c.�v���F��w.5P/��.��T�R֨��m�K�3�}��3�LJ)���4�=�V�B��.g%�]��!!<
^�*�}�����nj?�+Y%�d��3`]�@
��Ž0t�_4�J�I,�Vo0�D��쵈���d���jA7���p��L�o�m��ުԟg{u~����p�o�IbT��`����5�s־����}���ɘ����F�N�^��؎��t�����t�Y�x��XC$/����V� %O�9y�C_&2J�Z.K��;��QJ���Z�c�B�#��c'�V��#2.��#�[�s"�'�4r���\��w�^�=���6S�;o�ks*�Js����O�l�e�1������$C�<;��c���0�D8Q�["��Xo���B�����L&�au�D�f�=ڔX�)6oe�^{�c|�L����cVc?��y�z7;�l�����J��2h�_ү���4A�R��щ`SG��mۥ@�<L9�h	:P����U&:X�f�[p9W�+��}Ї�E����*ܺ�v�BZ�z��mY��G!-+��v�_0�uظ�(�,?�A��uF�U��	@E�J�Ć��pVDG��*�$��X�����aha����n��X{ˇ��c���ST�*;��,\+��Uɋ���������ӯ���p>�W��g3:ik���|bFR�|��R�k(�'���b�7�_��>��	�"�9����q�3���Ԃ/�M��U��٧�������m����׵�Q�6��b�= �6�(�"�H������p�y�ZÁ��_�����O�)��jI173-�ҽ%���g�-[*!� ���{zk�w=xrk)K��P����K!�5�9�R�C�G+�u���d/݅��+V��2el�9[�5�r��x�&-��m,R�eR� ^���'�}W��5�N��χ�l����F�.)��g�;�%�L9^���p��0\�M�n�.�k�cT���%�O�;��^%DL�5��,���)7�e6�����hlK�Vfx~V�E����	��(��G�<Ě^;�qk�Z쀂ǫ��4�Z&�_~��ΊD>f��[sP{��~�y��-P|�<�����O��ao儫#p~>vN�����5d�T���'1�P�9��~�\DM.�r�v�vV�LE��伈r�X�V%(8�@�ˣ���kL\�Ag��Ce~�R�Ͻ��XL�p���@��u�!}RzG˩�k0G0)Y�d!�]Tr�:>J����HoB,��'6EqFBߌ��j������yK2��?�w%�><$${��+i����6VK���Q�J�	�j��7�S?d�tJ3T0��B�Cʨ��YI8��鑳.��j>�P�9s~7��t�p��g$C��vX`�7�|7�j����:mI�o�#�'@�XۄG��:%SE��b�S"������Y��u6ۀ�.%�[�W�������|�����*�D�k��P�r�IY��śAɆ�$�6�$�!�L��\�$�ح*�Z!eK�b�)t8�j�Ƈ?�b5�5O�vH�&�X�zb��������۾g���;:��������,+'(�t��º� ��M�{���s{7;�~�>fN�u�9{R���C�8�m?�'�xY����3\�����_vA�j�I�b�����&Jy�#v�v�����{�g'm�
H �mX��V���r抲� �yv����P����f���1�A�JJ���9�Ya�3)�f	�����r��4pS^E�j�Y.������p�2�^�l���+�)�$_��YW��$98����r��	wn� �D������I�͖�~8�]b��0E�b<U�&}�-7�G ڱ��]��I��t�\�ElL?a����p�@r2n8��H-j+A�ˌ�^���
U�^����m�����N�{�S�eᕏˏ�`�/.@�b�%6��x�`�b��j�vfga�X�����ި������vh�z�G�W���I��/2�B��#�x�Tja�N)�	����9f�9��5�������c����NȞ���tI�5	]�mUB�Ω�
�����4��B�l6��-_G�����Ԡ&�j~]d���}���s��r��Z�ҕH�Y�c����E�hۛ��s  �Ӗ��SC1����ݓQ���`�����o3��y3.�O}2�3g"5��r�HSP������;�I㡜���_�5���"��{,�D�� �[Z��Y�-���縝&;n�Bk5�̜����L"S,P�{�HS[X����8�j4sZH�`:P))�@'�3��N�l_sB���~�<2<�'&������qa'�5�nO}9�<T�R뤻�{����b�\Z
E�c�#
�_�^G��И�Q
�w���u=����]'�hb�H�0څ3R���)%���z�1�o{��Z�s�n����ԍ���o�����j/ңNrw�ˢjUpX���/Q�1��L���c����z{n�5mS-�;��J�/B�9;!G[UU+���8�)����5�lkz9
gKfN�A6��8J�[l1���ӥ��l�J�j�������!@qz�b{)!���_����|� I��~3b��g�҆����3z���hY�x�q�N�9��<���N��$ $����>a^!������Rj��l�U=Z�S��j� �V��&�*Z����׃�����x��ê�@@l`�j�kI�$J�h/i��v-��h�R_T�U!	!C��$6��#n�?�qt�|�1����m\Ai.�������Ɩ�Ԧ'�Q�Ԑ�D��u���Wh��sg��>�	ζ�3+���C���,����Lk?����x�8;�����73n���z�cq'�6��)ָ���}��(�v��V���6d,���U���b ���%bMQ�E+�L4)%�m�VԴ�l=RD(}����7Rl�}��^�Wp?m��XJj7�����*�'��Z�y!�ocH�;���� �#�m?f^ΖFwZ����Y��nva�U��X"��֤h'J����n�J�� m̫�$@>G���k����I�o_�j1U�܀F����c�
D�V��S��U�M��3��GG�IZ�*)u�#�m�1�R[�d�˄��!,���&��s4YEH���\��m���ΏSR!�$1�a$���/'6U����`�6�k[	�V������l���m[0pbm7��r
<F-eB#��vR��~wu�f��>��r�6Y�5��Qf��<����<��]+�"��K��Ϣ��iUN7O1�SԾ!�^�ʤaX�A���'�F(�k�Es��F2ǚ��w���)-�ZĤ�cS�����2r�iw�\ЄJ�G�ԙ׼홼�`f�&��p����dV�"t�A�}�(��E�R�(�P~�	�h�l�xEÖU�%�~l7{^n݂t�h&( RA����L.��[Yd��ݠ���jqdl�_d�OW���x  -$�p��ߊۘ���ĭ�ͷ�G�2��\�|u��K�m�� = 4���w�iJ>�nz�aU�((2�kՠ� g
ԫ��?��l���4�t&���aBX��E��5����I ��Y�K52Ò�s�	��l��t�d'h������F)֤uǟ@��;2�=�7֖���w�Q�:pY�_�/M�0�3�8m��)�lvە����%�/��?~�`�FCa6u޼dO���,b�dC�%=����!��8DT��*a�$)�%����c������=ן�#����Mb�"���	EՍd�PlK�.�n���]h��\}�tA��z��"�"y��*���g�%y��c*�)���UPU���&Ֆ��nF"l��K�PV#���XQ�m%�xj~n���6J�X1�n�ݹ�7`����{��la@�_Ύ�DX���>o i�UwA�B0h�Lŀ{M�YF�F�rsi\�b�A@����Nڥ9�N\ �� � H�Њ#�;3I�_��Ěz��l(���>Lh@�l���C�lݑ�a�>�����h4��z��؈�	�la ʎ�'WːR��Ƌ���F)�*��G�Џ��yS��|�L�k�%3+R)'3�P�g*��ݹ塃�#C6���Ӿ V:���,r3��D��)A{<�+�<��Mf.8#��S�}�>�6{M���ǛN�Ɩ�*��·uB�N������4���T��x*�3��:�K��Y�f5�v��c7[9�����^��dY�(t��G����`�Di��&�9���"�~�3 C�{=�IJ�8\�/X�����h���W_�@c5�bp����x�֑u�b����e�֤>�U<�׀�l��{o�o[�7��Q���3�H޿����ٕ��6���*ژ���Gf�=�,U���r�Z=�õ�[y���L�SH���O��|aȋ699ry������P�Z��.l�뱛͉�K�2�%V��m�l��fX_Y��}��ـ���t���4�^�����yN����sA��=�,�X<�h�]gsw�Z���\�
5��-*�)ˆ���렠&$�r9��ć���R �K9Μ�e��5���r����pc�$ ���1��h�L���Z��)(����e����,�vP��Xhj�X[S����%Z�pr�/̙M�흼K���b�V �o殎�*6�0�������R�'++���c�����u�����ݡ�����50$�F���\��oٙU��YN�w�����؈���:pm�Rgjt{�T�$ac���f���}�&���_b��f��L�zؑ^O���)$��뷓�t���{�`.d�6ۧ�.��M�-ol��˽}��Jl��z�3�s�V����QB������Ir����e��:)!j����@�G�d4\���AQՀ
���L��D�&���8��ߧO V��5��4�&`�Z���I[�ո�IY3O�����i�C6\�汉�x�����L?��V^��-��͖=��`e=bl��kBA��P]m+�1�.߉RJ"e󫉚r�$��@���MčM�,x��mƨ���r��,f����@/B�/Y�r��I=�m���O���LLR��]H�Q�.���&��G��1Ρ9y�ǋ�q[¾�o�
G狃��Hq�����)2��b��̖A�bX���˝�����Q�ĥ��3���z�W]�Ӆ�7��ȣ�!��:�Q��߱MhY}1��FE�$�ьj���z>)۸�1�����e|��7�yp��Y��ΰ��QI��"P�j����dokt�?�l\��n��'\j�/��}�l֞`�i}]���cxl�>�pH[�t���鍹��s�o��,��hw��2�2�뭊��{���Xft0vEAd[g ����0����vg�@���n'�j�#�@:ؒ�nt��Sw�����>�/�9�n�Ӳ�Ԡs֭��F{=c�����b�o3��^5��s]Mһy�a�,�m �_uA�g������x�^��R��3g��;?R�����
��G�$[��b4�v��?P�7�CPm���TQ-�6���Oɔ�{�vvBR�v�Z8�3 ��������n�٤����5WY�4��u�Q{���{��C���t�_�$_{�.��f���>�n�:�g���0��_{�R%����%�)��x��*;\�2x�򗗦B�5`�J3��7��nX-�F�{����œ��M�p�����7��g��{�۴Jc׬���ǐ�Ђg���d��7��J����H�~3d~�֌q���CZ\�'��G��0˷Q�Y���:@��K�
���V��r�][M�F��/,3�p�Σ��4�~��&�h��	��{��l���d]�4�̅Hj7����_�dw��X�-m{����������<9�a�Ǩ�ƨ^��12�����A2ŔP:ju�<,���H�A(��~��&|��"����2�%�Uoi�z��&gk�_�w�6��1��Z��+�|W�Z.~��KfݘXD�&����@=���f�͜���Ҹ���Q�a��24�֓(�ꖫs!�"'ڵ��S�n�|ԩ����T��#�QK��6w�_؎�:o-�f!р�HHu?�
�oyRII�I"`F�#��Xg'e�U�2�2������*nn�2r���K�B/9Hz�M|n���bm#������0�T�g��&����1�����X���~S��oh�4k�ƩpM1����=�,�g����|�ľ�3&��7�3��Xzu�e��t��ю�뫷���˭ٚ}�L��}�bI!ǈV�f�/�IP�V�o��Mo�97���(2�E��Y�r�� G)�����z�^�FKy�V�ʶV=b`'� ����}]�]Oi��� ��J��E��tSN�gzE��FM�n�^%�J��."g~�?����Z4�BҒn��^֚�Uj�ٮJ�H�<Pf��a�M %��]�C:&��:88�;��y^�Ѝ��M�n��q!غ�
�'��,�o&�؆&w;�es@Z���Z��w��q�MSOE�x+��[��#���Wݰ��~?s���һ�U��,T��r�6�!����y~�PD�J���:K�6̶�����@W�]v�5�'/�p��E�
T�ZK�o���fk����t�l�m	�t!�6�z0u�-}N���T���
��ռ��;˧�o4)O���?�BhC ���>�a?��!��7~�?���.�|�j���q��"S%T��*���7�c��̀�R��>�H����$��zM�4��c�^���P{�Ś�;xyv�X����9�6`��`����
_��`%|���/_��er�]�3U���<����	:8�p�^�1,j��,B"�sr<��?������i�۰�EL:��Cn�x��4�d�˭��j���Ȝ�8J�6|�.�t��p��DB�l� ��cܿ>���n�f�S���-�1部B*`�ʐ�=~+�|��Ib8*n�����i� ���>\��83��7�������U\}n�O��Ԅ��2�R����]ͩ�ND�}]�][��L<������3���rq��[����M��$Z�^l]��PM$���ь��*�ŕ�i$�&���b�-F��m�U�8�.k�^,�hg�6�d�Rm]e֍U�5[�W�>�Vs��pe�&��U�i}Z�?�h(.�+-EqH��D>�����;�W۹�;��~�H_�<�[tǋ�,P`�
�P��h��ttҕظ��#^6�8Z��rMO\��6ʜU�T�\�L������U����V�/c�F7���R��>��D�$���ud?��;���k�_��,��_�����iv����zޝ��@܊B�2�H����8����UovbS*B�c3C]:1��V��GmW>ϒ�M�*�~~�� s}7GlCUX��Z`���붨F�0�О̜���YٲKs�y��:9H����K³hF�����9�Zf�ܛ���>��~��"�ݐB$�wfK�5-�z��C�\�H��ޛ+�v}�� ܦ-�g����9!]�I��6P�߻~G*&���n�I�;־�`�` W7L���6|����]��-}�fSu����`��h+X;/��w��!2���S�ysݡQ��bwi�l���y�ʓ�lu�8�Й��l�?tJ�+m�!�i3�bȔ��D�^2<Ӥ���u�585������y>�m)����B���$������^�X-���4�U��]A3��:W�0��
n��
V쿁�ul�A�d#-b�[WK�5[Qɹ|CU�$kp*�t��LI�5�c������~ kg���+�,]�`�ͻ�洼�'~둼�B�V6��f ڔ�Fz�S�*�C{��(�%w<�d�,�f�o�taHQD5�S�w���ر7ʏAL"���f��~^迟�)E�+h�5� �/]�i�5h�����HQ�4ERD����u��0�Q�V�֚q�P��g���t� ���s�y�m,p��Y���Ĝ�*�Y�$D��ɟq�#��0��ۮ��Հ�R�h��J�/�*�%V6����u��h�L%bآ$���{�� ��=��cԗ�՞���/Z���#�pn����ҭ�ZYqnH�⡆ۇ�>A4���bQ�1F�a��Jf4~�z��/���`��.����F�I�LJk�k��s�5�����`6��K��?�,��Av����'<xo\���p��t�SWÇ/^���l����t`;���{B��@���ʕ��P/>;��.��%����E����0�yso�~=��榾|EL�cz4Ar�D�+;�2��`�.���(��xs��F�4{t��s�����kq{��]��;��y~��`NC��cD�%Ǌ.���-m/�9�l��2��]2~�z��X�{�1j-	!�z�{�TE�o��	6q��a��\�m����Ë������]^�?���o�*<k�l�f] ��o)�"�S3��9~Q"iΞ8����as��A��\f���-᠌��ѵ���XK����ھC~�����{���>���{�8�R�tg4���1�4M���p�"��:�l�OW��7W9�&Z	N���h^�8����0�}>!x�/��O����ya�r}����W=mAl�m@k���Vo!Q0r��S�R[�u�%5vu��b�i$�s�j�8�����r�bo|f�؊���f�>j��D���}��ޞ�n�n��������V�[��KQˋ�;;C2M��y@�������r��~�/7���2T�[f���=_\ԁ>����9v��7�݈��ȵ�AE��ɼ��Xf�Q �7�dt	��:�����9����,�.�bכ����!ֵf�L�,��=.�����%����g�e�J���i���#��qqӏ'Nƕ�C�:�A�M�+��m{�t�� V��W�ee��U��'*h��$K=������es.T�%j^%{TvE�\��_��}����Ф�������E'>�)�U���w�I_{VOO_�졐����*t�#�����Y��=UM�K����V���
C��<¾�'�N��K���rH���AAW�����`�:jrIv����K�J��qxx�	F�������WNd
,1����L�bW{f
��#>�oM�.CGŨ%��|�s���b@v[�f��,Kd����%f�=pթ�Y-��\��~ �D�Ӽ�-�r��bPI��P���2��|�OrqY��drI�uY��!1���a@���nW�:���4���ӒΫ8ì�Z*叏"���S��s��FaV�<'������z��L����9yXM:�c�V����8;�B~﫺�����+�{\!4�?$�=i����y��i�!&w���h#�����)�v�@!�fJX�1�k;v
�Z�ǟ�� ���1�P)vZ�
�VETR��c	~�@�/G�q,����POy����t��jݗ�*�c+�	~߭�e:�V�U�`��á�"�W=�+OF����s苤a�;��`�G�L$��X��@��+o����}��-�B�	'!�r���k��"˚��q�?'�9����+�a��&���<LG�׃�!��^���^�{J	�?Uh�k��/�v�_��f���~�q���r�Q�3c)`�qk�:c�d�*bAD��Pe,A����`������G�-��ߨ7�qgH��Dbb���Uȣ�=%}T����B�aĶb��N��((֩@�����Ԟ����6��c��l�r��t��X�=g%#��E��X�NJ|D:ю�V����8pZ�M�9
�}��2���uWE�%�h�k1-*��hݭ��%P ?��l]D������dl���'������_fl�u%X\M3c�.��׻v�m�j������W�~�x��_i){��Q����1z�ÇU�dHF��t�����)(W�UL����MU��j�a�X�k�>��H�7+'̶X��o��7���%Zi�l���S�*\g��3�����5�����R�����b����UO���C,�}�����u0v`>'�2�����x$�l4�W}5년��(kդ����r��z1��)�F䱕8GoE�h��H-�D�$����/32�T��ʿ4=vzS���Ď���c�}q����r���<&Q���d�f�y8i�{��!p��*HÓa�`ͣ�K� ɏ9�JI;��� KL�7&O�)[ ���Lt���\��:�y��)����Yo�J������|��VJ�Y�����=`���ս��p�ޮ�%�?�[�x�mߦe��,��/ic���Vs�H�hk��H���F5�=Bϳ'Az��BM$�iV�z�as��T҃��_?%k�޶�����J�'ʷ��bY�l��c[|������ѩ1_A�U�tX	#՟��U�����Y}�c�q�����[�_!�o��N����;��t���/(��,�1I��&�,l
�U�05�UU'FuH#��+�ɋ��m��76�ZmbJ�]��?)l�bP3�A�H5r�i�['�Ŭ����r���J%ק��z{#8-��t��MN3
C�Ũ���ĩQ��}pFƇ���[�v��fZ���,�56EŲZ������GhͰg�SdtJ�*	ah]>�HG�D��Y�]����K��s�����^Ƚ�n^�}�m�����o��m��p�̜�S{|�n�z�v�����u�\x��|R0B1���F�D�С1���
�h�z��B2��-Q�/�'~,E2��vp��H]�
Jʫ��#bT��4 �����m���$�
��Ĭ)�Ȯר�Kߦ�F�<�@���9���7I�Wr�Y �M�G6 Oφ=��F�I�$c�e� ~�<�N���P]ͅ\J�	�	�+{�1�G0��x�����EU�������I���
��AŢ���W�$�Ok�R�K��\���/y��cb���@��x���3����ɗ�zQ�Y�7{̈�nH�����M]�����W���� ��-�j��8��".x���ʠ��f�e�k�-n-,R��xpn ުq6�;J��} �V���YR�6���۳����u���B�)�e1��#%�����=��8��E�XԊV[|ݍG)iuLqF�t�tZ[���y}Veq9��T/��ЉYDll4�W���Rbb�=K�P]�����ǔ)�i�ߡ���3/���GT�o�!at�yG����7�mz~����J���1�!S�m��ʍ[�Ü
^�o$�M8�Y��j�F01��$<�С��ō�(���w{��CE5�׈I�J�;<G
h2�-D����$8�o�5�"(LQ?FŬY3��;"�#�8�e���J:�+{�ۺ[x���^����S�_��~���_w[9n�[�Cفk+{QWY�H���r�A��a�;�)�}�m\�v�WK�^�*T�Ì_4�<�Ry4Þ�4g3I2�~�+~̥��׃�`Y�kT;K19���w�/�3.�����O2 [�oF"3I�_�oG�}�|���&��ߟd�>��yJ�!�<�̅r(�S��M�ْ���R��
��ˀ&�'�)����;�D�Q�'b��S��Zꎲ���%��7�MVop�^������S�eߦd�mJ���͋S�[����<O
&�������8W��q�[w��/���Hii ��"t)�ȥ�`;>D{���f׽ҡ�i|(f�݄p�&fn�L��A�|�^R�\~Q��`���I/�E����r�v�~cyk׏��ZlS��B���8��=��я}�*dZv���)�w��+j�A����{Q~k��:gg�.��ӓS��7E��M�0�4�Tbh:�:��2�{���c���ʱ�4���/���ɇ �e�ט������Je���$G�yMS3ݎ�53�Y��"s��x�� n`�����}��6�e`�N�Hdw�[��/����4I(.��h����x�w���f$��4�\j'԰P°�G]6d����}H�\��GU&���ΛR<��T蟛~��@�K΢Keh���n���6;�������w����/�?�:�?�*�?"�ԈK��:fٯ�tLqr����r#6�9]o�@�7x�7/P��OD����41�Zs��8�C�����-#p�q3a9�]2��׆f���5���k�R��M�Z�����|�n!�����%ֿ�ǥ�����0��x����a�c�7!sk�?z�m�b�.�sД��h�f_ea'��;}���5���7�u�=��Ҧ�B��g*~e��c	D֡,�^D"�rP��+Mk���J��+X��Q]�wu<s{@�YJ��E�'�o����;����vޝ+����g8w�Rc��h��O�҂'�����&�0�a�_��="����M�������3N�i
)�σw�|�� ~�c�z��̭7Mur����93W8SRXJN-���Qc��ykRv�N����_�K�~�$�<H2e�xf�*�ٓ�2'�F_�bY��q�ĸ�����<4��j�lK��V��m=ic1T���v���.w�a�B;��Ҭ<f��W�m�4�q� 26�Y�@��TӴ��� �O�C��J� �'b<Lo�W���g�(��t>�,qow)�VWz+N%�����Cv������@�KM'i������V��:�g�,(�tn�M�<{#u�<��E�bE�1U��}i�KS�����o�.�մ6��6�Q�i��j+9���������0<��OKm.��[:���#B�!S�>;�~�cM�Z�=n]�s,��5#�z���u���ڋ�h�!Ȑ��/U#o�,m����Q�Q�!U��H`������U�1��Y8S@����XBf;sk�G��W��a��V3<?^	�L�	�����ʘ�؆���Q[�U@�`7�>�D��H�~b�+uv�$���G�l��5�A�1֯C�;(pi����+6N�ĉ=�)�I����Ҳf�t<��d�N��Q���C��W�󋸫p� �m������~9GҲ9h���GP����������tr����Rǟn�:���6�;�1'9�^�K"����ȣ��������ā���ο�K�у�3������T����Py�r�} �%��й@�L^Fd�!�a��O@�v6�@�G��������!]p~2�^_�)�y|�YItc:[���5����Q>�"�i�͟�u���saq����>	��Ešf�+/�/ҦVL����羭�<��e�k�]�,�M���bJ�}.�z��5���R��򭯥G���.\n�A�
@��Ζ����e�&���[��2#%�,�j��Nju��n��:����Z�HI��=j��vm獀���Θ����d:���Vo��d����K���W�}I��Ց���3$w08�J�,��A���¤c���E.ߵ/�'������3h�D(c$��zܭ<�N�P��{�{GJa����Qi��}y�Rvu�V�.�O(��v�ӓ�ae'lke��{�C�0 ���\w_�x�l(���ə���:�]��8y�'V���<�1r �N�kK\p�O��3f��{EǓs��t����R��a{�$����E{l�}L��a��(+�r�~EF��E9k���?��NC��ƴtzuc�r;M�x(���p˨뽊<OK`�R�Er���	���Ev<vm�N�BX��%�����s���l�E6]d�\.�!�	�h"�h58'���>h���>']���Έ�F�%���MIz{�xY��f?Jx$���k]��Uv%c
��Ļ.�a�Zq^1�Sr��$�ܹ/ya��~���m�i�0ĺ q�te�iu�٬�(�?�������T���:��V7���������f��	�������|:��:���:f��R�hx%m�ι�v�^����ws��p�˶JN_����9��G*�k�$�Wܤ�@H��4W!,t���XEz0.���� ��{(V�-R$���JѮ!-x����D���g���n&/x��(�Qr��#r*��Z��,�+�'�>I��u�bv}�5��09n6m���6�=�,��l�KjY���mz_�*�+~�S1�w�]�����^�N���}�����Q��ʶjm�9ؼf5{��ۇ�GK�Ɣ��<��"�@߭W�S�/<�
�O[��s�����'�=�|��|��\����^�������o�S������·ǟ6�ܽ�V�ѐ[o�:�>?źrӆ�׻���Ԛ����s��)�7��^�jR����տ�I;��~�O�U@�S�����/.��1���_��N4O��f���ռFf��㽖���V%�n�2+�I*�sά]rA�:�*����;����)NѢW*��Ŀ����7'W:��h��3WV��*������̽�}\�FO��zU�+�޵���EM$o�]�7��p:쇦i��Ň�?\�������&��������υgrʴ��ï��,���n����;����}:���`G���}�����b��]�y�*��Ӿ�}�䜲~�����<ysm��e�o�����<V�hC�������3۫���O��ŷ���U<��۹�����*�ߟ|O�N^��n�m�K�zE���t�C����7v�u?���~���A��j���_w���=�u��[��tm�.���Y���[39��=�}�.�w����]������]�g��7'e������{?���s�����H��[SmE6��GqD104� S'���� �t���A�e+��#7��&1E]�Q����m��uW0x����sJh PK   �n'YXs�銙 � /   images/cf59327f-2b20-4f20-97ad-1ec426c5b43a.pngl�T�m�6<Cw�t�Hݠ�(�(�H�H�HK�tww*#Hw)=4���>�s�k��Z,��c�s���M���2>5  �WUQ� З  �\,�'�~��oh.r�����/�E8�gl' �������.�C*WE}W]GKW����l]>�;}�u�l��� �
��=3�=<���1���/�U�Qq��hZ���DĊ2d��s>�u>EYẼ�SP����L�H:���pt� ;�y�o���P(C ���ȁ��e�$���)Й%vݚ �������f< �٭�=���:*�������0J��	���� Ԙ *@F��u��}$�)IzFf�Y�	��$��;��8d�+9������%F��-լ�u���{إk�o]s���W[�Zx��d�Y�9��$����ʹ��R����a�%燷[�2S������x�9�w;2z6,���2���� H���m�z�#�2"(���	�X�w� �/�q�լi<hk��.��\�X��$O�߉��s�g(�4'eh�j�w����Pښ�ᣔ��'�K�sI�NY7?ι�X^��2����D����/�<2��|�|���F��i�ŅƮ����5�H�Y+u�7	з\��NC�/�����dJ���:�^� z71���'"��gl�n$�n;{��h�t����u��va�"��bEie*�S�c�#m�t${F�滬�k�уQ�9��v��@�MW&~�[��l��Kl7��v�^ݧC�>-x5����n���,��XQ,�����Od:/z�γ��Z���Ol[��k�c�,.&�� �U��"���mކW�L�x0
�����w���MZ��P�0��-R) U2o�Ng�����dt40�R�r<�:��qݦ��L�,%]�+�ä��SvxA�mc��}��O�C�Φ�U�$�b>3�\t4 (gn���'`{�'7|�K��h
`h�F��[Q$*��4����@����d���55�y���=��$��n��NmgD�85f����!oc���_ز� 9L��)�)��1��G������ڈ�x�N��m�0e��/�-Ħ��T1ɝ˟p^"���� ²hHF.>M�<�n��C�#�d��YT������sۅSV�Zx�������fwD�ԼX�n������4z9���|�����e�2�hC�~L��c��Z�¢}�Ο�7o%�ð绡�p��}�v�=3�M���� v3o@�R��:�i�'^"������e)��u�����_�J2��R�d8��'�s:*�U[kj���_h>��gr����͛<K�>sN1	H�=0Y�r���{����$�^e`�E��"d4,�S	?��� x>{�_;�˚ě��������X�J��T2A�@�'�K�P$��Y���e�R�l�MR�$R�㺪B= ���o��EZ��8K��`�$�40���Cˊ@1\�Y�ӿ���'��-��e�Y{����Cv�:�m�V��o����mj��Ԑh>qz�'!j(�KO����gn4��JyC3�M��?��"��`��M}\����{�\{t\S.j�3Sst�߫��/�8T���3G����6�gj6����O�0�=�EЏP�A�v�#I�����>�����e�|��}�N	��¿���#��+ ��RY������/��W���K��\,����u�>�u�mUx�N��&�n���K�*ޙ{�L�e]]�˹���M���Jюt�+��^<y_e�<�[2{�8����@��AbZ�k٠<�:��V\����A������/�5EGg1c}	��=���%��~�ߍR��p�f/i~"�T�>�O��:�� tw��f�A/9�۽�d3K�X����mh
���_aߒ���;��^��˻1$~ZJ���}�rz�=p�e��w��/q��)�G��ބ��[�u��](�l��g��w^�8���tA��I
je���R,.t#�o�b+��ڔ�7����u��H<�I'�g�����(��Z~Nv�5��h]�1F�R�Ç�pw�$sC�6$K��q������t�ܭ��:Uq�-�AQ����?Ni5E��|�o�ڭ�5 �Ǩɿ睳���3ﵠ��� �ݓ��Aj�s�>��t�v;��\�����;�d��J֮�����P�8�-�{���Yz�OMGi��Z�������O�'�{�Ute�P@b��fO�C̷y�8c@���:�������M�G�X���6dտk\E�j����l�dʛʴ�/e@��0����o��8N��
���]x�)���5���!p~�i����-3���Р/8�r����>}m�#�4�1��A܍	;�0�-�M��a���%�� G�<����6��`ȏ5مt��u�WtF��{vhb�Ѝ10�h��	��A0� F,����4r�@;�Z��"ŎI�]�[e6�ޟ.�.�v�v����x}R<�_�)2���Ǒ~���ms!"�(>p��:g;������(��E�n*�����c�ͽ�k�mD���3Z��&��s^���p�e��d^�36,�sl[��S�8��U�+��_����EC������?r�٫�3�Lf��,m41��[��@��a��偳�/T�N���H0�F��v�6��8_�)"c�J+H�ǋ�;�u��@XƣF���������������i��$�ͧ.�<E��FbH��Y�t#�I��C����XJ�Ya�a60��p�:��޾�B���Ft�G�\��~_q��4�~�_Y�rt�/�D�8$��Y&d(�e��)z�po�sqA���/w"���/,�ܝrWC[X|8�����9p�LT�������O��7_�8��vd7�����~zN��+���E!�V�F��_���r��m�m{_&�z����˄�F�7;��+t��i��K��
�>`Xei^K������'N�Yh�W�D�&"��ٌ��yQ4%� �G$�K�?�yw}G9h	d1e�����-�<�:n0�x�;?���@������\ڶ�~B���l7���[A��ޫ'��g��љU~�B��㭊Ac~x����z���,ɼ	D�%m��廓��j"�x;X��|��4������]q�{fY'��;�,h��fe{�[��(!����L�b�=EϬ��δȏ��۫G@�Ԙ4�KJ=�9n<ߵ���hu\��uG;�d�/]�-�)W��NqB�E����d�]Ha#�?J��c�F��zZ ?�]���c,���VL"zlO�1*�&~mMݫK9Qw����S�K뎿�_I~r�g�c���m��)z��D�6֝������M�b�0���.�q�5�ܑ_��O5�>𩫅�'o"kE�]�q|�u׾����s��"3Wz���Dv�#N��G&qz/څ�U���P -+�k#���7=���Omݚ���%X�m̭��`�f[��̋�X�#|�!�������j�H:�j� ���$��9���2����l�8�#{VQ���$����I�Id:ȊI�.��)�����?����d30Naպ� �C�
���;:p,��׫�$`�13������SL��׈�j��[�Ƶ���wz���y/~X,�2v%Ae�[s�=�Bs�ܦQ�7�f�v�w�
���p=ח�N$b��+`ǹ��B2�;�،�ƛᲱ2S⋢����S�[�%���T�d����0�װo����>��}�b�w�t���4��F��kw��@�Ad�}�<��cmΖ�seʈ��O�w�\ľn����%eR��KLli� �5�C0	k5L�����I� �����A��i,茽YS|<�,L����e�hX��Tx�.�Rqd:��ғ��t��4�E����K
���ʀ���
b����AF.v��FV� ��Ewz}j�i��T�sz2Q��,c�QEY�e������lG�E}%���Oz� ��!���$_C���Q���ǃ�O��r?����1��6��W����u؇��L�����;u��zco69\h=���1)��}}�!�\׺m�28s�fVes����RNb+��>R����U�ǉ��'�4~ :*	*ޚ�+gϥ���S~v�$��-�Z?��O^�{�,��B]��@JC�����(�:�ެ�/V4-~�`I��9��c��
���ײ����X�k@� �m��q{&]�
�����Lp��_�KJ8�9�)tc�Ke�ےϔkl� �w&���d�UZ��I|��)H0Q��A��Zry>���ˊ˽�y1H���|�T�g�<����[�Xe�>mC���~�~ؕ��sz�������E+56Џ#\���L�X�>��d���o���/����E@Q��Wid�-� qt�n�y��+����X.mԚ��yҲ�d��l��B���]S"�&? }�䑑�M�޵�^��ؖwU�e,���h>b�?\�!���Ҍ��e���N1mqz^b�J��.��+D'j��(����n�(�O�[��;W�}����r��А�+����U��xI����������Q��9��[_�[�x����RUi���./��^��N��1=��~��;(݅Y�:Etl���(���� �̠1 �|$<80$K]j�ݰ6|`��x��L�)	o�td�<��P�{5OA�g��ݜ��72�,>�H�2Gz�x��k�2C+�/7�`��|�^p�fvڕ�l�3bVr���<]m�ø�W� ~GNV��z�#���"��LΜZ����1&gI��O���L~�j[��c.�e?�
��kMS��G�)�<e6နO�V�W���C�D��qL��E���ic��䯗����{�n>������˕H?�
��	�/�	�̽���3�i���:8{<��B[m9���=&YI�,�B��iz��<�=	���X�l����� �	�f8��1Dߔ�zޥ8M��T͔��tߤ������Kk�o��i��䳸���r���l?`� �5|��G�y#���*�i>ɒ�?}�'�N���2���֙���I����γ�兛dmB���ӟ�c��f-�<����'�[d�fzX��|B�����ϙw5�@v�c�~u�z�c��L�F�~�rd2\���d}��"�����9:}�I/w���)���L� �0@5c���z�.yϟ�c3od�N嫮��u�d=d6�囗��a�v����!�w�ܞ�)1s�u1�2�Ѥ��@�id�T�6�%i�Ef���ﴞ�U_d�k.��>Q$rz���gؽ��S�SQ���u��>��.6��1WvsKnsK9!��dZ�_��/e��$�wC�|��
�(��y�f�e9ܲ.:��l[�V��~�㸄V�IH�vvn��[~�/S���jyСl �jf��y�2>(�=�����&H\��%���{��t��	=�8��G֝�WP0?����/ ���o����d����ߋ9��\:��7�c�H^6x@�!;[?���v|�RC��1��R�& k�S�ud/�'3m����($U�L�'�Yh�����lCx�xƛ�֐���Q&\��U��TG�!-�5i���X��O��o<�B�u-�%�O:�C(�S��v�"{���͗���B݃W��W�)��?{���!��u5���>��7��dG]�r)b!+�AQ��>3q��VO����2!cPϕFv2�즪Ө(p���ӂ;v��/���S+�����J��?�0�Qj�u��xF�Q�R�c����HA:|�u�J�u����'Qe��7Ue�;"D�nL�f~4�M�5�1��l���2CX0��ݰb����E_�l��9��L��A˰��k�� �Ar����uzG�ӳ5��aQ 2��/t�j��5p�LF�i��YD�;�N
 �5chŏ�x>G'�hQ�9�L��uK�u���&���Y�t��[�f,J�M|�X��S�)9�;߄ĦD���C�Ԡ����a��y[�%��v���*�p)W�D�f�Q���a.XM4ף���{D�O@"V���Q;���������}��^��ɪO��hf)�gG��_��Nۋ�%��+��Tq�;?�c��'.��т~-��W��T�05)OpYփt�
L^��\�\mw�@���'k�Y���8�߄�Ғpy��A�R��*G�|M�h`�,�l5<����	�	h��/�Kr��"��A'�W������x���$N^,��0���؝�i����Xr�w=���*���Or[s��{�>;tI���E0��?�7��9j�R�p�)O=�f�U^�B&,��D°]w���O�tz�/�AoE�=<��d�%������+�Zд4����~�Q;I��
"�DM,�����أf������p�U�+�/\�L�^q���eGY���N��/qh�cKHwmC2%']�L�:0�Fe��f9��	 �&t���0o	�����)tZ�4�K�]�<���K�t���	c���߬�3F��K�(�<��%�bՖ�#J�齷%�@*���>�� ��#$�􆼝��&%���1���)&i��Z��`+w5��:ݍ���*f��ѿ�d�|?3,Ji�b���<^T����p�ņk��0�|����ۡ��܋S�W�>}>�y��+���v�#Ba�h�0��,�0�q��)�[�l���Dis$�)$>��7|�o*�X���?|9Gf?W]�ovmmJ��'ZW�HJ�bC�xٶ��\ \cNU<t�L���Z:ª���+��6k���v	�j�[����� K*5�`���	h�U7��S��]���1�o /���6kf��U9�J�;��Ӣ� o��`�>���4Ma�hd�`�_���2���\�Z�����ϸ���*^�]?lӎ��$�-�h��R�u�H�r����� ������bv�?�WU-�nV���d���w�T5�\JH���]XL徂����('��5ֈ�z���jjK�Y����Cr�����V1�rE����|)mR��4�m!	W����j{Z Bui(5w��lg���5뺂V~����8���k����#�ꜻUGe�U ��=}���+�U��q�`l��)��k���r�g4�ŕ��M��N�����5�E�1-�	%H0���'��Ƴ�A�{�9�C�����nf�,���cm2U��yI���c
.�T������7��F��R��3�u˪�d�h��ڋ�υ%Ju��}$S���D�	�&���,286X�5#G�q�>4)?{Q��.�ۋЎ8
�	>����:�] �̬�q�owZ�:�u��-�m݈8��� ������D�ñ��Ñz]i��l�"�[��?������k$��S׾���:�k"�
��w����& 	"T��
��۔�$T�h4/15�Z�Q���Fl�K��!An��ݷP~6���TPp�E9�W[ـVT�F��'|(��n��3ռL�e��}��짢�Ds��SK&��m��(�	t�j:ۦ"��.�m��aU�x�d�\��^.�����_�w�ӓ�dS�g/Cj`���_LB�:�m�F3�pd�M�C�����i��o>�Db��J��d�+B4N
��]&�;�ߠ�1C������z��.���l*3\���'8h�Ǒ)A���l)T��E0mT�᳑���;e���5:����N껫Wo�Yr}�����s9\6�>dj�T�xfd��^�=9��;��[��x��ONQ���E�3i�k�x�9�l���[e��O�4hl�e�_�QST�҄�����+�"�2n�j�F᎑�$��T��j���e�Q�"�H��wl����~so ���+����4׏�:���ʦ+�缬2k� d�M Bm�,�ΦMq��a��W��}B���BkM�;����;x��B_�㻢�>u��D�7�������ז�`Rk�H-)R��y�#N��	;sUFt�ө�6�$��Ƙ(X�葚�@����[����Y$m��Z�oK9?^�lgdOk� ǂ�
7?2StF4�[���n�pv����Ҷa�с�y�q#R+�)6�t+k>x�ѧ��ϰ�zQ���h8�55�sf1Qvk�v8�K�D�%�%!�.�G���|�HO,'����o��k�1��Ntdj�c�2@QY��S���^d��5�AH���a)W:/3�������P����=D����PK�G��CF��J�yk.��f��a�N�>�<H��(�z��8�!��M��vD���4Ř�Q6��Ӹ�	 (ԏ�Ea���������s	��"Ζ����!9N�q���)@���T����l]��i�;����u׹�K����ƺ]�>��7���e��^6�,ҷm]{
w��(�[���J2`���A>,����-%Rd}��.�G����QSP�R\�Ʀ}��E���y�)��)�ζ����֩����D~vO�[G�m7���<���a���H1���������q��������佌0�rdP�`m����c�e�O-����b��:�x�o]��C��ĻDs�$\Z+T��ij��;J=#F(����+%�(Mtej����o�U���e���"�%6q�C�F��q�L�__ѳ�y,[�o C~b�O��b��q��5̤��B���1:ZU�����|Ij�1&��xlj樝f��y\k��Ñ$�ʄ$��XQA}���گh��3��_����D��!h{h�zYO��l_����9P��m\�R0�F�y@�.!_.�k=]j��>8%�%�,]Ğ� ���+/Σ���̜�5����r��uL��r ��7Sc��:��0~T�p,L4�r�еSW�b�S�=#���Mô-��D�}�eؽy{@in����F������|��W��@TG�j�ͭ�9}܉���q�<�8����`�?X~-�q��U����%�D�39+�x��Rb��-^�:>�������;
"PყK!˻ER�5M)�r���l<�YD��w����p݁OZ).��A���S��s�D�Ɋ��ЁK!�␍*O-���s�{Ƚ����w�s0�s�kB�!&pfh����I'A%�1Z2�Or�\�]��j4�j�������-y%�%�o�K�b�H�}7\,��7����̡�M*F8������>�fM	y3]��'�zry9ǎ��sP���ђ�#�<��A���J�N��'Th����Wna������s���jѽ������9�))����l6�/!�m2D�mM��f�%F�d�#�O��ZoE�WQ;q\BP���u�t���)����l�z�7�ެ�)/-�s� �^�hH �����6�h�W�\Tյ~HS6��Y�ktl)��1l�z�������I�E�h~�5���殜;�;����i�衴3;�r�`υa�1 ��R���$A�[�%e}�fMQ)՝���hǉ۽��t��B���[�t�x/��
�����u�y��d� XU�n���H��S_,>jۥ|�?>@/������խg`�F�8�dy�2���_�bd��Q*2�xn:ۢ�d:���|�ޥ��L|��R1C9���9���;B}�l-.0�y������q�/d#�ц���4��o0���Tr��'B�����~2Nt�=1�[�a�Ù�bCx�[,>�M�lٱA67���,���oxĞ/����Db}��}�;����,}=u�_Q<`��|h���?����^r�3'���'����W��d#��o��
�}�`�,5D#��`�u����2�)9��SͧW��*���sJ�!�0sɈ���#Պ�1<6�]�
�I�p��0-EJ>kF=�f�;}��EaZK�����׀f�ʞ�8�_���'�hY��c.Ð��8�w���6~XUg��}(�I��#����r����c�fvM�Ͱi,�S��l�PH��������ټ�,�X�3|��D$��8��7��T�-��yBb�/"C�?�W�+f��T	�����T�0˻�^�1]S����`�Uf���l��a�w��+M�>!�g�e_nG���B*��H�G���d�>��/muZ�/�K��/
�̒�b O�y�[��,W�rkX��uT�B���S�.t�ĭ�3^5ݟB��@��J� S ���UM��7W������6�;aT?~@l8U�odK|�����! M/]�����^��u�~V��M�Gp%���}�����|�(�GTsJ��٩-�nV#����Ա����	�*�E�]Fng��"Œ�p�⮌Z0�C�V�qAj�Z|8d��viRSf�+;�r�������a�8i%��i)�qf&��H t�P����TL�$j��m�ޜ��w��Hf|Q46�V�f!5(뼕��c'nl�V���$^�`�^'�]���ۖ�X?'�W�E���q�[���-EtV�q	����J�H��/b�,v�p����3��=�!����hi�VU�4Ŵ��A��۹\��ɲ�F�E �+��06�C��#�H�1���up��p��L��|FaM�}�+�S�����,5Z�������="��ň�"��~K1[��9j�c䠥���i�Q�a��<_�7ft�8,�|�5~��њ���g�h�F>YvI���ѡ�왅�&����#�	�1j����J�xn��������-�=��J����=A�P�;�p�u)e�5Z�[�`���@�Ծ?��H��/��Fg�}��.�MM����{��?d����&�D;AF���o���^j_���e�$��Bs�띩
SA* /�e9b�J�P�����ԚY��iT�]n����|ᥦ$�d���?.�4\��M�PsE�
��E�(Q6���aE,�������u����`yd�
���e��7
�c�`��>a@x9$*L��_��w"��i�sؓ�஫�@�]��+�p�|A��'���Ռ�8aHfX`���|�H�W��/��n.{&cX��]�X�`�N\k��vB(K�D��I�ģ�n�"�zeͭ�A͖E�k9�We��d\���7�%uh`�dp`�}����k���Ԅ�X��/�U��~0�m�z�E���'��Lϛi.�O��S��t�w��J[=;ks#pSi1�����Q[�^! $8��������+�/*��ʼ�Vu��H��U�F�gK��軠5���5,]����}T:���+��%_���;��-�n~_���WO����^���j�1&R�G��#�.W	 W�YdQ��)�[�c��&��B��|M��*RO ���1��#��y��l�j�e;Y����%v�@������w��!�	�hc���d9�+m�-�TW�x�zkR���E΢j�5(U�5�|i�DOy³q��6�QID�v�6꒿�h��!�M�T�,���l����*��sd��_��X�bJ�ٝ�)�vQ���`cf�M�}���Q�/�d8�+)�/]���hfi�zox�Ϥ�c,ą�]L�`A��&���|��5i+m�_��o���א�qZ�������J�����>w�I6��ؐ
1t�=O�l���������ۀ��Q��3IJ#�ӽ��\k�b����rRϲF����fλviȌp��gt���I�.E���!^���"�zt
�����g�w��@G��v#6q�V>������Iߍ{^��Δ�<����h��yŠM!������(Q��E}("�z�����L��q�lJ��'"�v0"G���gm�+�pC���;�jTx��G�N���}l�Y��w��2�0�;��RF�����;f6�S�G|����ٗ
��^�� ?y�̈<&����r��y���e2�U$���U_���4�*�
,xH ')_��N-� dՀ^��vg�����!]���=66K���]���A��n|�9т�R��	=p�8'Ѳޫt��W��jp��u�d*g�Qh�M��*d��42�n����쓌���
-��ܿ4�>
�"OIȆujp��/�+���@�eJ$?.����u�n��J?P����z�͚΋�ss�o���T���ٞ���k�����ބH|���4Þ�h�,�#��ynL�q��A�`E�A䛵ܪDUשZ�8#Y�z��O9��+d�N}3:�R�p�|y�O��G[۶�����<�B^>:��dxБ3�����HW���S�<|�^���<�-F]�SϨm������"Co9�����]���g�'!C����X�����o��=�AQ&^A���8�ޥ��}�pN{��Vo�� r��@I�c!���br��䬛K�6�H�cb@�NS>�?cոx}}�уh�]Z�vGk����^�)lk6w���!�5��2Ic�99w�u�@rU+�g)�< � ����fGu$dH��_#�Մ[��OP	��`�g$���?�Na�r�ƿ	of_d�bVu �M�:�lK�aKbMy��V��0U$ ��f]�¢ϡ��p�@���6!�V�>/1 
O!;u����?�vV�A�P��']pz+th	��5o��B��l�P�ސ��58{�=醻[1��(}���!l�@����cY�3k�	Q*�KK?��1�d�&`�g���F8���)��?���KP1� {��MR2���bIz���/�"+�ُY�����^�M�[Fo�{�AQ6�(�oi���e��B?��o>I���*)��.H��aΑ{(�=$BP�8**
����޹�ɖ!ݯ5��@�9�>}���}��,�X�y#��.qz�̧�OE���jI^��}?���x�Jb�Q���@�Q��Ĥy����Luj��?����NG����\��r�$1E���"�O"4:�>���'�q���k��C��z*�l�2S�����>*Sǐ�i��-]o/��$NE3ػ��7Ф�+5��2l�x�jy��EF��4�;܂D~�vf�W���呺K�ٚ!P	���H�A��U}į��G0�K*=��}k���$�x��V�y�KN���=�)�����X���%�5���;f�c�o����J����¿��z�N�����k�g9H�!��R�/��KqU]�3b��w&��Z����Р���X��d˿���s��Qo8.h�9�o�֩��"�!�}����k�v5��1d|ωEW�W����E�	q�!����l�ŀ�=�_��u�%�":��dh�������B%������Ym��>�/I�̀n�ݔ���4i	���+0����D�'*@�����%���gL,m��8��
����d�����t�f����į�cüe��	U;�إۀǲ~A���v
Kjդ��ɕF�G�F7f�ҏ�	a9D&��W��͑��@�O��+.5N#-����n᡼#�gQι��;iR&����9+���*#00y[~7�����<�)^��k�ޮ������d	W#�Ҭ���*�>�\�n h5}����i��m�|���Aؠ?�F�G��� ;���8ݲn���-˥����,U�,��w�����dj9���aai�P�N�&��2MC�������,E�����NxlA��HH�>�5[[)pz��)����w��m���g�4���&���%����eŞ��g&-t��6���������"�P���Ba|�D�'7N*0Ա���/��}���"�:r�Zo����^�a�
�@�E.]���ہ�ޏ g�}��^�M�O�����˹k���8fi�ܲ�O�5kY
�э�/�Y��F?<;(�դs�!�J����'�/q�:c-�>�:[?i�6i˯v�8t>�'��gs���Dn� �&��s��ڐY�k�|	����5�I��9�ɶ.;��,Ňo�S:�5-�뗹8].�goO��,�����^�<�ey��ړ����~�]���eYh�t��n���hj���/_��ez�9!��s7�A3�μ��{\���4��g�7R�xU��6k��\��V _���,�4SP���`�yȒ�b�\T:�K�W<�nI�IHD�3Y~r����ca힋�}(����TV������t
���~�P�P}�u���oa�W�O�ϰ t�<|�����5%?�5������%���}�M�k=�P�����m�+2��������i"�^�./V�'���؛���o��;�_��4�H������f����:�1�["�k1��X�{�s]_
�e�ۧ;AL'm.�$LN�I�[Am.QBK,i���mwҬՐ}��9�����M^��ꓜ�(t���}l�3 D�A���� �i�Ub��j�����}������ĝ��-c ����p�N�D�<����3<Zj:~���sϏ��?���E6Ndڎf��N��x)OK��4����7�k�o,�f�ŇG��"�ӿ��$w��	u��0.���}�Ԁ�q�����F��'�N��@Eb:+���](�������+�h�o
Y��Y��9���is�h�5|������k��NtR���ᡫ���^p�ʖ�*g���r` Ï��l��Td�ڈ� �` ڳWI����9
�(e������_�%��β�i_�����l���ƙn)#���`���
�|�#�!Ig�5���N�e��ޘ��qM�N�p�=$F���_j��2o_�M�/p���y�SFi�wԈ���u�q�c�ј�A�p;ӀR�S2pl�+L%@�:��.f�l#�����鮀�( ��iC�-��}��B5S������1%�ʲ�[�t1�`}|��q�WI��Y-3n�oI�hڿG�m��$R�kʪF������>?;�w�����sx*���%�(�u'��I%���S�R_�B*����{��4O�%ݘFmo-K��?�&���?���\-��-j���;�)��q)2E
RPh$:���:�Az���>���M4]��#�3(!֛�a���L�ՔH�V/�lu��y��bn�1�l��sS��\|��ac�{����\��c��1�RΆSU�uS�_��8蓎��r�)�A~�.�{��<�tn�}8�M*v>�T���P��<D%��s���](�:��̍�W�궰'D��ʢ���v{��SGT�#��Sm�EC�p�2 ���|.�B�w�(��Բ�)Sa�툩1R�/j�kQ��NF5Q h-#.N���� ��UE�U/��Kc�A7N�Ys'�
Ǖ����>�A�?�C�J��(DpL}��uʭ�t�;C�=6f1ss���$r\���wZW���(裒C|!���zm�I��v�F��y�dK5a�tiC�� ��Y�ﻹ�	;�rj�#�2[Jf�a�#$�ȧC&z�����o%hొsq0�{��/T��'.���~D������J�A<��a���?}��{�������<쉂�Ee�`y�*��-�e[9�b/M���߼۩n
}\��a%��OD�借V-{Euh�.UI��
� �6�R�<9w������H8c�,f����ɡg�3âUS-'�ZhpD��N��b~��!|��'�UZ��b��NQ�*�Cs���ΰ&B�*�ks, ��%oo6����a��M�ڣ��r��qc'�lgCRT��K�Ñ�v�"��?��S�d��X
 0?=����%J�#�g��a�y���'�!4򌋏w�uK�#^w����?fVFl+�,��H�J�^��.;G\ۂ�~�n�%y��@�y+>K2��{�ZX��m��`:�[1����樦�V��S)��w�����t]?�G^l����~�NS��S��sM�a$G���F��푢�pF}`M���t�[�Nٱ��k�Ț?b���BK"_a���ڡ�����|�s#i`�&.no
�~�4� j��"]_.zI�]`}��|���2���a~�h]�z�A���c��W��8�	ׯ$��T�F&���L�� ��V(�q�Q��Ӡ�`�?�&���f	��(^_d/lXe$�~���#q��>�h-Rd�ޠ�Q�R��<��5A����NYc�Gx)���V�O@���A�w1T�Ǟ*����.������߱�i_?�-3T��PD_�NU�������V������AfL��H�v���Xib�5 ���h,fۣo3"��bzFz^Ѡm�`9�	�"��Zؖ:{-�o��������G��&�BU�TƱ��ܷ͠}Õ�������d:��/�*�\neW���eL^�ĭmh�Jq��/�s{D�Hiz��v*<A��_W%v �A���ϐ�B3�j&D���;V�y��7�A���)�?P���/��|NtX��6u����
6l#���(�:��g��qX���ͯ�T�]�5�d��ύAQ�\� �Z4,sm��=��Ab7��R��j%�1�J���/�1���mAX��z��k?���t�F%_�'6�W��8�"��w���O9���ޞ�e�v{�����au^*͢���&��f�K���?1ahs�����렠ka[v������GJ��������2["S�/S����ݫJ�[L�����d��T]�ȭ�WU�0j���0�f�Z�'�H�lnņ\�����V^/1y�U�r�� [�%K'A��C,<�伥4�ew�c�U�k��A�7q��Z��䯷���T�c�V�y�
��.�;�h��#�P�J��I�4�z�܁�� ����qQ}���0�t#!ݠ�t���H#�Hw��4�]�4Jw�4 � �����}��f�ٱֳ�z����l�[{p���lek�!�_8����ym���Bq���,�"��vr�M�Q�|�U���Od�h\ҧ��Ӣ�̳7�*5�;dP����:�v׹�|od�|n�ž�e$�~�"�1�qw���H��>��j�#��J�s�E'��~T%}H/���56�/�=��2�����wL�_'}墄��C�F�ۨ�I�@���[�w��q��Nb���[��麱s���H�z���p��/{��&��P�09��Nx?[���J�6�� )�$O��#K=�M�C3P�r/�n��:�ov7��cc�n��CD��u��v�0�^>)��gm�&Ŧ�=��0�/��u���4�7���^����#����!�6U�،"k�DC5�8�8����I�s����^ƀ��-ػ�7V�zfxt�}#S����r�����=���ů�DSz�D.ũB]T���Z|Ư����Q����^R*��ׯ������������(��ӎ�3���\ˠ�r��MK����2�N��Z��>>�c����߆���l��~3 ��p%֩k�o*�s89���&��A
�̆6&E��f�s8���F�J<gvҫ20���;|u�Ə�����k[�$��8[�u��'��:܎���З�Tpq�o)��}'B��u4�8**}�#��b�����u)�����a�bG��u�t��Ѱ���B�7��mS~>�B�+��g���@:��j��f��=���ɋ�'���>_N|b|�Q�f6�V�R���9T������g�8u�f��u�t��o����'O�j�s,��q����jvJ��%���O�{?4M���W�k������n��f�Ƞ��}:�o*�?�b&s�)��0)�/����� �}�o���H,�o�Mi��Gj*(C����u#�|���qGQ��rb��E��:;��۟�'�juY���)��h�������'eN?�gw1L��-LE���E�ZVð�%����A�8K��1����b!%S3��+Q�ݔ ��:�ηmd�7��"l-���ty4���������Js�B��Sx��abj���djQ,��F�Ij���f�$Ks��P��~K��_�`�F��>wI4�����x��|���Xϛ�@�]}Ru%p�e0STTo��pC[�5���׫B+~������eyK�vrC��n��B���L7�m�z�E�[)�WAx~rQ8�b ӿ���}pHb�ѽ����(~���o�#?s�s�_����X4��8�x�A�3SS'(��(`{(��y$D��o�\������]Д�t�#k���+�Le!�}����V=������J52�J�p���"Ou�w�~�S�W�q&'K�(�܂����j
{u:q��+ݪ���?��f�=R�tN�b&%��<;�������쩮䣇�/i�|�٠Y�`,BV�S�\��4/����@�J�o�7&vr`�m_�[Tebϣ�#㊜�����B��Zm(���p�)c���P�L1"����o���4��{�c8��N舀���&��h�4��T��������
]ϳ�{?�H_-50����">��.��&�U�%���� V�.�A1������F��.8 �W�f+�� !�u��j��^�R���eښ1�CB��zDf�}�F�7����}�_#�h����(�?���,��u�W�)���?Û�i��ȁ�%��B����{X�
Y�kʝ����M	�*_�I�g"'C�WWX�
%H5���i�D��PɳP��dfs=[�v#�Q���V Gn�u$�ß�@�I@V߁� �B��t�C�V@�n��xN4�j�}�w��o�;�K� 쌖����L�uqr�^6}�sqX���u�C�8s⿴������Ž���d��N��}�V�v/0��]Q��!fX�8TB��y5	]��ytl]m���L$˳��_���v7}��A1\�MX��Np�SNNƹ]&�>Q�|�@i����L�cZ�qSTY4)�Q4��3|�5��ϛ���}�'����r�l��o��\���ڻ�ϡ�	젳WFS~�\a�Ls�#�q�ab.��DcVAe<�q��-��%I���,Y�z(��m΍<�wC��~v�˃ H���|�a�b��,�����|�D���"��=	g����_1�z�����ag�k�X�cI�q�w�����w���e2Ɵ��CP�.Pܗ���R:�:�] ػ��9g��lh�^���uݞ�����xξ�Yld*��5�$Y���%Q�p�����G����־� �%0Yy����P���_��#��d7��!e�["��<6/�����Q��A���~Z<��V�2,&��d���!�����}E���'���s̢EN���Ƥ���t �D\؈�n�8y���"d���>[�l��2TJ����T�c7����_��=�d���Ol����z\t�g�e�]�R�� F�E�{E����GZ�w�����*�%�qˌ��9�T}����9^������aR6᫠�Px�3|ZW�]¼�d��6���lзtx����[]��2�G��q���w�
���}�8��8M�	�:��Cs(Z�����J���������\�=͟�m��.�$(���|9�Y�8��yv"��$m��H�w�Tn��E~y�~�5w��~cGC�<.[k>�ٻhh��~D�h��'����T���K7�Wj3]~]��9���hr�W�D�kc�=|K#x:��S��N����,�Ԣ)����Z]��T�6�b�XҮz~�S��z�_�z0�P<�"ˍu���t��q�+T��HϾX�77+�ǿ����M�8��s��p���_]�=x����!j_��rr��/�fq�s�"MՋ8��:�A� 1���#��jƼBA.aj>���p�[;?�����B�y��
Yc|o�oWv��JH�	�����p@�*�����?�}p��?F�N��?U	 ģ
���13�w(�7�\�|�{I\}o��s�a��{?��9ϲTW�
:`{�d����b[�f�"�NN�{2���t�'5������;8�^�����iT�8�O����b����;����Yׯ;�9%�Xy�̫�GY�wa�����O�Tg�q������X�t����{�!X3�N����yyעZ^�Q���9H��R�ٍof64�
�&�T�ä�}N�q.���o�t��E�P��j˓a����n��6]:����yN|�f5�z���[u��[*�F�c��"����Otǳ�g�8��gOi݀W|���
�������:�<���&4����X��EV��!c��������R-�V��U����������e���1g.q����N�S;�uRW�nu����E�Tz�R�+�7Xܴ�����'���L�(xE�n��&���3�C/inGJ�A�����(��P�RGGez�~�60^ͭ��Q�[t.ѭ�b����Y�!�8B��r����	h:*���q݅�v��*�*Ǐ�)���j|��Fyu�9𯚼XDt<��ф�+���}�%��񚚍"��Η���;i����a"�i��O���ʹ�w���*��H�1~�ڬ�[Q���,�`l`s��"P<"ݲ�'�Uϲ�����FPβ�d��[���Λ1��Ie��^�O��o���]��/m�Rn� C� �����i��d�&���K��`,!��۝~ߕ���_x�7�D�s��Z�\�>�?��mj6]���贍|���ﺁ�̣�`����^p��{��q��s�IX�c�����!�ѿ#�˵�n��L���m�l�������j�ύ�K��� }���?w�f�(���� U�������F��IՇo;>z�/�jG
��eW�"�(�ē�+Ƿq�1�+,��-��{�v	��Ff��C����a��U�p��P���O3�2V	]���"��F�~Ss��?�x�?����䒛;�6��.L��ݡ1�f�*���*膾���oL}X�28PK�s���0?o�+�`�������d�K��XY������Cz!��8�������A<�nX���@=����*�kab�N=FW���3| Ō}�h�
]Y���>ɸ_?���S������b����V������Y��&x�˼���ۭ��u��ȏ �������Q��Ǭ�a�W��Bg7���s!�3��I�W�c�kc�8�+�Te<h�R�BcU��yd�Rfc}�c�$T�DK�4���l0i��g$�<]ot�G��*�.O}�x~�z5zo9D`�Ġ`�Y�5z���Vt��YԡÄn��Ir�M��1���t�����tZܮ�*���P
�������J�h����Uj���h�!��CL{�:^�C����gl���}��rSr9��N/N�i^HWc�RU�`�8T���龸��
PY���|T.d&7�a��.�΃oIÎ�3 �X4Pm�����>@�o7w�������$����,��.k?��`�Cl��AX�{�3�/l��ؤ��H��0���d-��xy��K����X<B/wް��7+ϧ!�sx/l�Y�L�����P���X'2���'���9�����JI��p�8��˻J��+D�pJ��A��Y=K2p�(��꠬�HX�I�#�[q��l�cܓ0@�?(D��E�П�����A��\Ā絥�����o���8�ź<߾O��c��}'���s�E��~V\�aɮ ��pd��7B���0E�P��O�;e!���'r@|�~����w�yQŏ�N��v4����I*h0>�4�
K?$�ȋ�Ր�eZ{�?$�;��9n2�(vDx�>����䭑f�s��t�`�Q�:Fq(������������d(���������	�cH��W����3)�X8_�7T�ܧ�,AIP� �:���j?a��� ���
`����S��I��"���)(����xe4��|����D$L�n��wn�Y%�����-|�i��\Ďވ�&�P<��`�[d~]{'�گ��1Y�"HY4xm��N�/h%ǁ�o/��.Y�㓲��,��L��Y���3G����Z�Z�2~0Alv��u�9�vlņ����`G8�G���zI6C�b�����{�K�?��Q�[qb��mz+�Ĭ)��?��aq/<�ä���X���I� �{g�h��z��Y�wD���V�w�g@��P})+�l�|a�l����� S��@p����uL�� �������"�뺁 �6��7�jN�K^c뀂W�f�Y��%Zl�2��R��jk��r����<��.I���*�-�Z�@y�d���I(�n{L�|d�8g%�[L����C܁�Ip�/T%Z���NM��2N8�K,�h<�W%��|u���I����â�E��;�/�,.�&�
L���S����t��.���@99q���̡��9�nIgN�Ӷ\�K�'h���kT:)�����#z���������?�g(����et���e[��O+�q����|�.d$�52A7�C�5�z�/�n10�����`���v[2�u�Gm�?W�uu\��E��"�+5��ÜBI�rK��~4���H*�)���J�W)E_نT��
�$�D��$�KF1���������m�))�xq 0~����ĭ���oC���z�* �>��(#i��i��,�~��.���p+��N��#���b2]�OL?�����ʍ�2����G�G_�o��]����mkB������m�%�4"�T[����u}-���YuR������9��
)഍}��[N�2�Mƀ�ˡ��~K�7lN|������7)Rh���Z��d�Ϟ�69cX��'+�)::8���'��y�We��*�������핀�j�Yν@�jYt5����Ǐ{*hG�f��EN:�Sn��ޗOQ}����;��;>1�#O[Ky�hR�G	�]�}T��d��v*�7G�y��z�BC�s�3!f�-�{)�xҏ�tL�@-��Q���bO�}n���.���~u��8������eaw�٧o�Y˾z�2\((����u���Q:*�4�4�y�ʴ�k@�ǲ��`:��q��R,�����I�n��ص������^�1��έ^�bd�
�I�2�~ms��Q�JYN!�Pe�ʋ��A?/>�;tT��S(?���t	5�����9	A�i⎫�(��Z��W�㠒�ā�Y&f��A�`�Ш�LM��P>/�j���qU�m�� �7E=ڭ�>�6C���i��2��=j՜�+�"d��vb�-�B�
i7�=���1�l@s�o>T�y*"e��Sr��!�wjf$%����O��Zu�#ֿu.G�Z�WYC|�|��%��C�����U
&�w���*��&Сe��tn��}�E��	��R:�-ɗ	*�yK���������'� �/Ǜr����L���#R
O�����e�˝��g�r����ٓ�T�W��'˕2����F�B3y#�ux&�M5(6q2��r����*���F�˂̡dn�d��3ˬ�6�� �����I�W�N�����0���M�h���5qr�M�:J�'���瓙�P�)�4{���=l�t1���&���Ԩ�H/�����/�]�,�������a5Gp�@�����j��zꢲf���G���� H�|H���ӛ�	�~2��5�ɺb�wn)��(��
#�륈�S.�6�>^��n���(u������kt+}��M���,>
����,(�{9��7�K�YW>����ײ�Z���):�)�W��q�5�L{�`Gw|F�X�E�<��yY���=�L"1����aR�m����a2J'�����Su�f�/a�=�c�-�q���{�� +7�_��.B5�7W��@]���G��ǡ@�O �ON�Ĥ����'����I�����9�V����C�Q�-�-� �������0�v
�Sֻ�q�����˪����J	��c�f�!�J�-N��`����v��I������&�1�'���
�M���{�{��]�o{Ȑ2� 
��N��E�Y��t$��x�N��<�A����M���/�ػ�L��>�ɑ!J�n:�--e�rm�3�O����C��y=H ���jdR�ϻM�9_���KMf�k��i���I3�V�p���r��p��D�ߡX�\Q4���kOYY�r࿝�bZ��F�lU�i�8����9;��.BU��[�$ w�42W�٪�&�+�s�J��#�X�������f�/��* �UC����Z,U�5>�1�w�n0^�O����[:*=M�5\h"m��J�e��++%��t���t1џ��d�\S�ȅ�
4�ԛ�`5Nb�G��LP5bw�������{	Ǜ Y�+���q��W>�ш�Ox��t���\�d&�.�ۦF�iab�dy.$��B&m#�*��q�b���3�2 Ќ��G7��AObȝ#(-X�3��hGt�UU=�n�r�ƀ�����_ޠ�ℨV>���v�ة�[J��)� �-�_˰7�q���F���L�2�r8��jd����3S#���	6�J)тC���?~����2���ڱ���W�ŕ�ߟ- �M�vQ�-�$�k"���dc���V�ˍP�q\7���a4g���ptk�8_KX��6_[�8e(1�/,ԙs�p�BB'�_��g��ǡ� ��c-��f	E�A�� �@q�t�&��6*f���vq�鏌�����lن���У3����{�A���
,�aG7�:�2�/|������Z��ZR9��C͋�����êO8�X�K<A���Fp������,�����5P��V+'���(O&�bNhP�d�6�@�o� �y6o�-��iD��"��{�-E��\r ���ع�FHe���O>|�טG2���s�D>_�u\�_��A�,^��n��ĵ!ff=���b����;ۮ� ��ۯ���P��Cž�WӮ�Jt�	�R[��e2�]�_����h�WU��6+B6}�<S):�m���J�2�?�>��A�ؙMp巣��D�)f��������&I�ר5}�h}Xnu����G��ߣ@.�(7x	�4���'��p�:t�_��q݀�4D�`ڕ�(����RW;d�̌�yX���hX�ZUP4����S��)ftY�4W�Q:��ר��z��"O٢��foo�����y̤c��
CW. �����!_
�+��j&����MΠo!ؖ%��Í;xE;�&3�>�Q�e�II���>Wi�Y\Q?��μcukS��es�wS���z-6��A�g/9�d��N8zd�~hٽ�xx��@���@�(�/��P* ���\���QWWd�(D���jХo���ػ��ms;�����A�����/�98t/�b3��Sy��E��jo� 05�AJ��l~���okuH������p*o�سﲜCc�1˹����ǿ#W3Ks	�"׳0ww�j9���&r�B���hݚ�D����Ԓ��C��"i{m���ˈsYlW��d�N4_�9��KqX,�x�49"B5����N_ʹE}�c�b� ~�#K��C�RU��w��
W!�x��p%=�9B<�a~��r�v0Z��29ۀ��ER����F����
�؃��4,���ߺ����kKx �ŧ�$H-@0ݎ��܈����=�����nFO�A���d���7\?j��y�
��8�̆��`�H��������M�@���m 0jd�@��	���� �����ueE|���ĝ@��!*C�H���'C���q�a󱽃l�V ��he�j�E��Y�*Gc)�.#�?X�O ����"J�R#�߶(�K���FT�/҉pOS�t#)K�T�����l�I'�WY7D��x�iC��M���>]!���P���z�1g��4y��!u2::࿍��<ko���`��l4��
I��d1�0Y�c�S��(�\�J���W@�@
3� ��'��^�k�PßX���X( 74����f��N'�ۍ5����L����:\LN�j��X�rYQ1>�^MJ��~�F/�֏P�L��kj��C2C��EA��m^5��q~���!����a����Z���ӕ��斥<SD-�f?�r�nZ�7��94]�B\:�2R��,k >3�!$T���@KX��3,���R��p�����0�m�:��fK��c�Y�����B��0�^��x#�!�!V�_��M7�|eQ}n�w;|5���kr�\�|�x��JAE�C�k	�C�:9d��Ԟ����I��x0�B �,���vÆ�sX?�Y�Y�v���O�f]����:=/l�x��:������;��V8E�S]�j6�W���y�̈�F,O���+�J���B��F����C������p�E�B]��$⢎K-�Bw�*j���I�YUJxK�����K�x�5����;���|�ߤ�M���ݜm?I��l��KԝCp�X��l���L�*@�����e�楎*�l���QPsl���_��;G2�'6C!�w�|i��շ�x؃��%6o~��MS|��m;�J(�D�H�!���B�m���W+�\�Tf��Amw��K�2��|�������"e�,VB���i=T�G�%�J	4b$���2���@�u�)�_�4��9t$�x��K�C�ZJ��+b��?w�pb����wI<-�*�	Ke�#;�U�]֡��	(0?2�a�i;W<j:�X���b�+�t���e(���i�GC`>�m�$z��<V�su���ܬ|�w�L �/|�>�6�&h�8:Ė��qP΃������1*���(�0cx��K$%���%s�N,��xHR0K���z��X@c%��O��LB:�%���(����f�>����Dbe-S��(y�?TN��!?� H��_��r�}$�Lg��B7��A�-�F�uW
���Ǩq�@;
̶�� G��j���W�&4s)r!�SiL��	a�M�U�k6C!�9�9�O�/#�ҫ1�Rś�{b_t����y�ʡ����C {�;?YTZ��Kc��!�	�/&�5�x��+���6�k' ��{���*B�Cr�ρw ����:C@4O����iI���yȎ�Js�"�c#�Ɏ��
��r˻����2�����M��_}�j�cP,�/�M�J�IH+�G\�\՗С�YF�R8_V@t���uE�O��eD<6��'x]+�d��,�&Yp�x+P�fN�̡��}�{�{����&$��,>�����ǋ(.C=J��|y�c�y�?�(��eu� W���4͑��	�<	9�����1i.����������_7t����uYZ�׋thG�}�&ȝ� i�RO�y,ܜ�����~��E��y�F�/,���K\�.�������Lڀ��A?VJ�W,P��ሴ���� Pk�T��uH�(&`���2h�cCH����w���(��N$�	F�������H"�n����2k�|=��u��j	�����fT^r����w_����%`�������P�WL�@m9f1��ͪ�G���m�u+��EE7�,�T0O�]�Z�v�`���i�~�|C )0b��!��0|�" �o�ʡN�R�,��aM�p:\�O�������p��\���$��q���1:�m3=_C��Vg�����  /9�'z=� �	�=_@
�0 $�]_�,*�6��eQX�K�^I��������dYol�:]�9��������8D��,~�G���3��S�ϊZ��q@|�0Q� ���}t���Q�����/m���r�uv%B�ri�>nB��� D�ģ�6ߢ�@N�o�s�f��MK]ث�#?��7*ʱ��y<���I�0��0��·�;�㆐�|� �����,��^@UC3U��4gn��K`�*��Y( ������y��x#1HtAUbAԔ�&�q�{m�8(<�{sH���5����a�ׯG	�D�e IUy�<�NP�q_�^���zZ
j��/�UV�[�٘L^,�윓)���3S�8>�Q���T|�0tEw�V>*nj
���iL�N}�2�ɿI�gL�����E4��	ȩ%,~�3(Z�bR��/��B;���X����\
c�͍�#��H/��?&��B���;�4.ĺא�`�,�s�!h���@���W�o����׾�c��Bѧ��F��C��Ƌ���ۼ�$K+uAo�}��įtA�#6;<!?������	���o�!���$�t�B�)w�'6��z��ɏ��R2`�UM�b,A0%�@������nҋ��>��Ht�r�NwԀh06q�:�r"�Y���)P��Yqk�\1����>��=�X����.D�����\v _��кɑݻ�]��
+�#.�pǛ�51S�u�S娴P"9%1��m����P'��&i� vv�Y�`C�R$ 'W.l,C���w,��hu�g�>��4RgpS��bu=�"�
�8[X��c�x+��ڸ��*Ǥ%fl�vK�* ��r_߉E�c�2����=��h���
��kni�'Y�'6�|/�&\x�����+��];i��}�|M䷧�aȑ�t�n\�=3��CX�.��� up��(<��:�@g���IigjP�ͳ�������ʟ`, ��	ts���8&��w.����K�a	ͬ����g��YGG�O$�p68����r��k���C�*=59��;��sL�c_c��e	��x8?/�����:[@��^�a�$ht��HS�cN�o�����#6�&�h'�\���?F�c#7a���}���n �{C��+���^�(�r�X ���h콻!��!���B6v󓞟��<svAy.���-Klդ���!��β�����O���p�{6{D>͗Υm��3�|���YAq��Ȣ�P�uD��i�Ħ^B�A��\��- �)�|�'Zl���uL����@���p�t8B�/n#�b��x�(M��r�YOd[��KS#��1���۳�i��ށ�-r,$%hw��Ԥ7!����F��Ua��G��~��S����!kEK-��!��B�-! ͆�X��RM�گT��l�; �h�`��ի��k�n��K�榧q�v*�ʰ��)S��W�W¥,�����ީ�|aw� q�sٰ��t� R<�e�V���yy�s��|P���5{
H?�����%V*�1-�U�JJi[��*M到�x��c�Θ�ʕ������|�x�'�S��o	�7���YM��s����kf��j� �H�]l�3��C��+�1�����j����������G-��}	L]��!���J�2��/"�6�KE|1W��ũ�G��"�-����%�3$V�G�.���-y��D	�y���CѦ7���xd4k �ۈ7t��w��
��+�G��(G-fi�/�f���@���H��G
� R2��h5��9 ��6P7P��Ѐo����m'~���W$$)�u��
�D�0vU�ý�9�yj�g�r�wO� )Eac�?�>�Xߑ��shf���
�K��J�u� �pM~f���j�'ɫB=rX�4�s"��u�|K�e�����k�S}�F$�+�����aE'f%e��y�'�S����4^<�\����t�|=��p�G�=q�"=���S�?զr"�E�IC�dq����9@�M�mUkO�ԹM뺕�B{���H�:�L��n�Ef���e�����_�5)	�F�d�?��C�gD,]��Ƕ6�tVw���[���6��������H�$�oX�r�qI`���ç.e�Ʋ挍-�w_9���;�^M�Lifa�/�i�#nRH�-����ѓ��A�[���J�^kC$�]�
=�7YWLUӘ�a��oe�b�\KE�h�l
��jV7��(gV~"n��Rn��W�H�ֶE
چ_2+)���Ij/��K���t���Y�\����Sg=���|�.���+�է.ٚZ�7k�0A/� -4�i�mV2,":_�������Ɗ��kf|�*qw1�y�:�r,��v��ݔ\��}�P����g)Hj�8y�6^�e�-f�9:��P�vR:����@����hQ �_ډ���4�Ц���Aj&ס?E�e�j"U�;џ����e^�`2��8�*b�Z˱�$V
���K[�C���!��>�ޤ �+7ܿ�Y!=�P1�:��{c`���ݭ�]}��[B5��H�v��ԇ�t_�D��@�lQJn��ŭ
��R�Z�����W�H���-���OVU�֡����BPU`d�|z����8(���0p!/��ͫ%��a�T��af�Ӹ���aW�����x
���ul	��l��&��z�7ӏ��*����k��%!Dk��|��b�v<o5��M���e%���}��|�&Q���>6��ئ���@zM���\�x�ݞ�9��(��,�ߦ��]e� wц^�D?o��c�v�Ґ��h�k"P/�7�v����������X��)�D��7��tm����U�˩�|Ǒg£�%V��T�}LT�xB Am��G�-�s�
t�:a!�$��N�Q5����c�$�c�a��'�3vx�_���͹e_�B&a���>�<߶ P;52+iL�ׅ�N�:�;�J�������%;��������ZNn�c=���3���i(�� ����� �E�{ns�K׿�Y(g=��3�|�X��;tK�ǡǪ��<ou1��ܟO"���][������l���G*X|��pZl����]���z��Xq�N�ٗ��%U�?ۨ��W(��ܨK�k�`~3��6�czI�f�?5�^�튮:�4�v��9`�h������{����C�d�g��+-�yB�\�N�`D-.�>�Q���D����TKKc�� d��H�Q��n��3�Tc��R�r��}���u��h��ݗ$�P���V���?�ڝ��w��ɭ�Y\��h����V}���������P��"�
<;pq�4�<�#s�G�~�U;xMqҁ����]޵X'��{�*�����5�f<&��ӳ�.�{D�ߕ-?��@�9���n�$<�<�4!(I$؄��XSS���<�	R��R��B����rX{×���9H��츊	�������{/��Gh�@M�T�cN�X|�@aߴ�����	��Z�{��L�?�0�O9�+{ɟ�Oph�)p	���h_�bj���2ϜȠyab���c�)S�L����+�SK��V�Ч����;������)��%�z���#��5_D�l{TWk�g�G�罉������e�.u�i)qKQ=h��3�.F�@c�Y�[t�O~J�R=���4\�=�~z�J�x���� �Ϊ!����֔�e+3o�˃�`��͍Q:��\�9�^��2 ҂j�vZ,h�(S�� :La**�>0�8�#�D�nn7SD���Ֆhq? ��,�&��,�����?A�W��,��K�i���km��n(�)�L��ğo�68�KP?��+�Lݨ#t�*�yv�d�3��d�oʫ��5�]���V|���(gbJ�!b����?�d�$��b�.�^�$�;��Moj���C���퓝 �pLr�r��%�3�6�L��� \��,�n5��h����]���>6�d#��%�>�3��+��W�;��O|j�R}�4��[.8�bO(rӺj����S[N��t��O�M*rs�ʖ'"��Y��[���%WSD(��uocqg�L��THP��ia$3���ֱ݃BI�n��H!^�㮓$HI����iP�$��sBx��{1����{ϛ������}��gR���k���7����ti����N�X�� v����3��@��������E$��e����Ԇ#zY��=
�8܏d���[
�?�D��mY&��dD��4��ob�ί����rHx��aC~ӯ|Sw�eq1�~Yg>��uMy��׾�,��lI/�6f�G���I�Gdw�����z^����w��mM�r��T74���u>�}�o��	���X����Z�9�SǪq���V  � �cj���;dqݕ�g����q�hA�K�`�\����i �Q�V�;�������04d�X]/��I9�x�ZK�w�	����&��@�k��$�>8���P���;�{��b���8����0��+B�.�`�<_�I��}�{�9O���7Y³�/�8A��u��)�p����2[�|ۛ�A�Vɒ)z�SL�<�;�� N�G(1rp`��8����Z_�jw��*Y4i'���Y3j:��/��$�-�#*�� ��M#��޿0��7��[����)��W)O�h2�|n~0�|��Q������R�^r1�~79�,g��O	�ykVL'��c�ύ%#A�	z0vF�Iix�392�κ��W�;M�d9���4fHX�x����Ɲ���L��9�q���F���v$CSO�+�����;3K�6X^O�v�ӷ���E�b��א��8�աc�OOlVϭI�,�	'C�5��߇J��2(���e�͞��:_�r��l؇�I�Qg��,�3 ]J=���
��UƏ<��xټ�f�IJ����R�d7��9ږ���h{��δ$�SdK��<�*�"�S"�A\�e򛂖/�3^ h��+:�6��#u�㾱�y��m#��V��Ұs��?mlsv �t>sQ�՚F�ޗX�/7�;�P�<>�w�	��e�&��H%{/������(��B�__X:��ಌ��0��xȕ$�cI����bJ�z����Ç3�k ?}�[�@΢P���fe�?�*�@���R�Gw�.e��RE@�(��f��9�S̻W1���}y�Y
Q�xp�:���:ڌ�_�m�'��_^�i����Ѫ!��n�[6��?�
��H�j4��5�?�� |����7,}�ʡ�ћ���E�or?<2�����SQ�=$	���.�cT{�{�~�X@Z��Q�)���E�-dO���X%��x�W��<���n0p�$7�c(?��c�����}`�M�_^���Y{ �ɲ�V����֔��V�c�[����%�]cM���7��U\^&rZ�><��X�$��V6~�k�m�{���I:L@f������V���	JC[[x��B9��7-�q)+����g��;�PƊ� l{3��^�yo���m�!��8�Ɵ|v<�4 ĭ(���*Wߑ�dnT��Lf���5��++.�����oR��:�þʢn���0l��[���͏�/V���w���6gx�m�	&��y�[����k���>�g��a�������D�1Ϊ�0�?�j��n�Qf�w3�ʮ��!2%Xէ$��2 N�$X,�����[G܍�W粆��#��o��J�ܶ��Fv�R6UE%�3��<����0e����m�y�U�Y���P���@�{�!{�z:N�@F�9g�H=����;�]���(<�����N�Ge4bQ�I�����5�/�H�ۘ��A��Q�h��@+�T��v��wE��f�5��-S(�`��r0����8�$J�%��!�*���S\M�5:�{pww�w��\�݂$�;�݃Kp�!��������?�V�S�JR3�{�����9ӃG=|� ��q� :�NǛ����Fc0�f��>$9#J_䪼� ����9�jғo�M[H[�L���>ETs��Q�~> l,-���/d` ����"�oкՂ�,4���#�>9~� �Ȩ��mк�6�ҶF{[��K[�/��G���ɭ��&+�N�E��yL#F��r���R݉'4��&�j���}iz���sił���3�G�. vѯ�?!�����Bf���Z��{W�����z���:Y�t���p7A����z�1�8�&ǩ��t{c
�U��g
���.16�0��Ve�����4wH ��#O~��u���F�k��ل?����p�g���1�՜�_$!_�?`���6���[-x��d�z�ST(��%^U�9�&�Lw��Q��1�����&�:*=����������WO��exPv�l��ޗ�CT���xs�op7򴞝�U����M�x�~�z1�����JXFދb�'����Z$�t�=�`]�}RwG/�;��>o-���)ԠyY{�]�LY���ވ�R=\�0ZKV�{mkί�o'�c$6"|YJG�V��[��Nb�L��B�sV�����˿5[7�E_�G�`B؟io�(���~n�;Ǥ� Y�'���~�Wѩ��֒u�R�|��i띔�D(h��C3��/O"D�A��ƀ�5�Q�PzS)�`��	�<��\!�K�p���^�m� �Sv��ń�^g�N:#F
�jy��;W�%�q���X8�&#G�@x�F֖ݟ�O�Xx�V~Ub$�h�z-I"�$?{}�x4qLˎY�IC���̪A�h��<���ѝ���	��q������i��2`B�h�1&ˎ�笖?u�*�E��!*�Bd���J�W%��ʬ���=����lR_��ڴd)��~{��!��u} ����S�ma7Tj�́<�F��d��l���IOJ̄����;�6�:��Q��,��S��Uo��<�6�~�	L�{J������UI�g˷�qId��_п�¼'��`)�����!�u�K5V<i�����m�!n�������J�ۛ:�(�.=_�G*8��E����rj<Z�5���6xr��iNѠt�SҪ�����&��~֪���{�F�P���Ni�Ռ�^�G���Y�ӪD��r�z!� ����D$8I��Q��mKY�N�-�B��ā�V��\$�<9�̫_��C-T�5�'�BYao�޻�͸}^��x�{Pw}�*}�t�T���N�L���Z�����E���*m�7�����ᤵN�)w&����{�}��;fU����6�%\��9\6�Dt���b����j-�.:�2�V��P�F������<g����)�A�!\����ϔN�\���`ժ뢥���4:�9��G����/JbD�cbH�&P��W���D	Ŗ���JJ�\�F�F�I��-Z����J��I�k f;�Mo��>!y�`���TLf�>'�94h�lP������E;��gT�"yf���J�z�/����)�N�du�7�����;�YFX~��R�҈���4&��nq��T!3smv&zf�����:ܾ>�lJ��JEc���<s\���<'�����H���xc�
s
�Tm��$X�0D��;���&�Vs��?��$%�lV:a&����>sb=��=z�D#�Yj:�d+�S�o�~���3��;�,C�"b
�]|x��e蒗���%�� EƂY���	>Y���a�e�Ņd�6����7�g�^#_�����t��m��[M�Q=���A��	zOe���4�V_T���3{�i��4wC��Z�"э@`_
�Y0�tur��?Y�<Y�֖g�L����zy9I$��/��F�9�����d����%lxNo�=����W�T�M�ǎ���h�1��@ҨR_��f	�61����y���=-�?�&��rV�h��*�K�:�,�^?|M2�mM�� �V9v��ѫ�*`Dr�������yz��Y.�Y�W��x�&��9�w�0K�ռ2\w�nH4q�Y��
$'����(Z�V�"QG��2Z�5Ԕ��O4Hw�x^��LZ��I\JRz$VR��:�����&���������]�����qfT�(��$H�Uڤ!rн7�A�X�Q�۷+�����Rj�đ��>��H~Z��e�`��<`X 9%�~��? ɾg*���S��H�*w]J�ND���I����'�m�)��A9ip��JL�h�Ĉ�����%>�y@@:�4/���r3@	���\+D�-�D[y��溉;���Ut�9Żp0ɵ��R�A�S��ʠY�����]k�ߍ���w��.�,Wä��g�ǚ{~=����Tۃ���h՜�>L1��.��B�l`$��5D~L��F �w��)]z�3/Q�����\��*
$2�n�*q5(�4S���|�2�Q���SX<���
@g�OU_������9�����G1o�wp�u�&iC}�ar�b���L�wT�1�Ñ���t��ް��c%O�~)���x�>����s�F%�*�uĹ�	��(���=��}I�MFy��Jͬ�A*�,W?�����-]��$��'�$�l���k �e]J�1�rVl��w ���a&f���ǃQ��d+Wĉ[�V�ɽ��:j_�������}���x�"���ϒa��F�48�Л�"Lv�6ō(!��������}-<��,�×������3&l
�j����OY��0��o枾�iYSY���hm����uѦ��G|�1�+�1�A��y���Gg.���,��N��=c�S4PP�1�3I�����ͥ蒡�]�r;� ��z̲�4�uF{�~Z*܀b�np�"P<'���'��R����e��	P��O8������W˃N뜺����ä���Q���_��m�7�#�lf|�&v	I�%����Z����)��N�!��sn�D�rS����Z,��"��:?�`j bh�k}RL��>��b�&������mj��sy���9�z,�"+�7���12,�K��-@�ϤM��Ҭ�
�bx�%�W� ��P.��4��=�؏��@I���Ь�x(-��眄[6��F2+����Q8����YaAlC�\�L\"�=/�w9���Ttdz�ɉN� ���Ҥ��4.{1J���'w=_���5E���Nw<!��f����G�k�j!���2ǒ
�Ӹ4Z�_(�]N��
 G��+QN���y�X�O�!�\�2V#5N&_�іo�0 |�NEl��Y��4�$��!�*��
�b	3�����P��G�v��_�!��͵tA���/�/�y���k^��:
%�T�J��.�h�z��Xڄ�#\�U�7�i�ʵ����J ��m@���U�e	���n�I��;���z�}*��s$�º�La)��� ���|ǩ�#@z:x��}�ϸcZ��LB�Z��iZ��2D̉�^L
hOd���b$�
����HU#����d�tW�.�4���ezسY���I:����S���ضke�(��a/���1oj�]XV��g-K�_ِ|���D*�Ts� G��f���Ӭ����_��'�֫#O�za���.�h�|)�0Qr�g�K��Yx�E�ӖVd;Y�s`�aRhA����AZ�c;ЮV�#eD�o�J�+�|zʨ��Ө����*�3*N����L��=���Բf�aY��نɋ����Z趣,�ɥ��OMȁZd��m���c����tBׯ�F��p����Y�q���z�(wV�O^���+���Xޣ0˖=��z��g���6>J֮`9��E�qU  M�E
?�I�2��yO�T���m���(� ��r`gk)�Y�H�j���ȳlB��^`q�y_��ih�-WCa�A�	�z�qav�*���qj��v�DS��Ng�h$�� F_��^��6���r1tvtY�	P�3�	�z8�{�
�ś�c�q���ì�(�\�=T\A��t��O�L��?�d���?R[�3@Ub��)��R<�S0�(����%�g���Y���IC*i�lד�Z�V�Q����5I͌U>}��9/4�#�l�c]jl�{��%34�P^�E��u�����cY�V���a%�ƃ?��8��'�RF�;Яi�^/º�m�zg]�Ty.h�sb#�J�Ԝ�w��d5�>��uka�O�I\�崂���ia�4]kζ�'t�%��A�r=���(mX�	�ș�o�0��7&��(սb[�� 8���0Å�o���|2��8w��=��)kD��I�ŋ�d�����I#+��ݽ��e�����k	�͏�@ar6U�a��x�ìv����iC�� _.;�9(n��Y�ʧp]��Οk�����6kPh�"���V���:/Z��i�km�G!P3XX�C+�{�Ї`ghh~�d9�
a��%�q���?NR%W���1;8���%��A�����W��������x�e�@�C(��k�a�+��+����d|F�f�LO����Pg7}���-��èF/�FF�_Ү����nis�9QY�f��M|��� ���Za��G{����4����y&C�kmM��4�gF�iZ̮�k�V�Ƌ��7��X�4�������	J#¿C�������1����:�Y�<��P�7��O9���׺I�9(C�0���vF��
��$�}�8y.�����3?3��٠,�ph�Y=-IrԳ�5Z2\�#���6����>�����{��#Ɏ_ln�@�R����h3�?���_��[l}�X$9�������o��=מJ(˔7^2�>m��/��ԿV"I|gv~/@z�? ��ME�b���h�"t��P<���`y����ꃊ�w���e��R.���ŷdmkd��  �&���.�	'
2�b���L�{ꌧ�Y���L�7�(�ZpX��%����p�������f!����a�����O�/�����8�h�ߘ�Ja�|�ʗʷ��s�t�f�܅j^X�)y������NHr�<h2�!�w�+b(LDG�%�{Y͔[��~�p�\�2_�:%�E��r�S��lQ7*zC�B�����&�^��G����q����0�Fz��7�F)w��0l�GY`���z�R�@_�M�0�S;�����5Kȣ:�òtK��;�h<0�Y�S,�U ��(�x��P�&W����>r�mVE�ᨖe��f�;_���Y�.1�����R1A���l���G���|�as���[���h|�(�ը��܇�\׎��s�sB�9�]�\bS�l0pWf{�}��"� dF{�G�]\���~�N��#c�����Q���e��*��z��w���D5uE��f]=�W���6�9Y{�jo@C�8����������)з�:jg΀U�;��٫�î�
���ӈ=F����$.� �Eq��[�������ˬ=��0<��O�&��-�׳��7��w�z<XI�������:�@�Cݠ\KO����:���b�g����QO��c�8=@1�Š�.�H�[["ӧ\�����Xq]\&��w��Zw��7U&�����^0�xK0�'<�c�g��0*T��,�9��ݛ�P�4Σ��"玺���(�"�'�f/0Ѽ��M�B��p4��<���iR�����
�a���ﰝ$%�Q��.4���*�3�H��/?�ԄI���5�y
<��!�֕�;F�4���D�,A��FK'B'��S-�������>�ǁ��韗�T+����t)=V�S(G]	ͮ��+���4p��֐nB�X������n}ģ�5�J�Y���$E�������}�4����D�t�Mo̪5.��o�	l+/m4�)�����*�o����Y��P�'��$dJ�M��	�e�jN�x9ܝ=�|�QB��zQa�˂LL������c1��O�����`H�-|Ș:���p5�������}(���V��<o���D��@�n�|l�ykRв�bz��[
��'ʹi�=I^I��HV��J�ne�9y'r4�ލT�D�D�h���a<p�[Zz��Me��Q����]��{�O:��NφEX��ʺ��Yǂ����Ig���N�T�'��?V��������=��0A�;I��!U�{���/�^�d���2��r��	[���<���G�U@�i�A_;s�EyrVh��k^K��x`�?����:JF�:P~m8��`0��u��d�/8�a�ۨS�&@㫞���F����7��r��d�^�bҴ�!�,�3V�	!�w�
U�B!SL9��p��`��a�����i|��]���v�ߛ�P7�%�B���d�ϐ���s�A�8�c=�Y��ň�]:ģ3/�&o��0,�|�5�_�x��1h���<��+j�؅͠�,o�-��B���cC2N�B,���%�)ȅ��p�����FOv�s�:G.���I\�phYH�f2v�0��D�W�l�V��Mq�`؏ߍ$�n�/�W��>i���	�ϫ���R�?z��؜�[/�gx��ġ�v*�:ѐ�Y�k!t��B����u���l˖�h�s�5b�F�J��*ҟ�i��g|��c��ײ��Z��h~�<�<�;�����1�[�m4T83�""�h�i�'�#�{GW;�����G:�+mZ V��T�����׻]3	��ĺTZ�N�2�d"F&T�S���1��� ���r���=c��xQ��d|��i�z��hGt��Hd���V�M���l�հ���������K��C�.c�C�T��0��Yy�6R.��$����&��Bs�D�Z_��"��ڐ��)3;廉o,PS���T =�	 'L�.�k�Ǧ��:��\t�v�V�Hg/G.��ځ�&/�h��� ����J����`xQ9�F++<�xc�{��懎{�ጓ�!���=��u�ߋ�����,�Gl���CM���L�m�5G���q�m����`�Ţ6�He1A�I�6U��@p �j��/��MV���G�c����N�1�h����)%��9�no�coR]���@�xR���\��j��}޳��rW#e8����z�W=o�6�Y'�����[`N��P�x~xI�����Y]-G:O�~u�_Lm�o�Xќ�b��������	���
����P2���������\3�<#S�Jj��d�EyC{ĊwW��'K���e������(��?���V ��/]]u��v��ygy]�'���O*����q;#Qv���'���]����d�v(���g f�>��"�[�ל��!��d�l1��d[e�&�OQ�
�g[Ggm��T�(����̹~��;��cf�GO���-8��a���w��(6����_,����R�<�P�a�<��d��Qn�=�@&3�G5+}�2�B�n��Fط� @凮\\��U��!1b	8CUd��Oa�|.<<8A��o���q�(��\�:\^��>$���|]��N��qSqq��#s}�PP�x.+�b|�~3G����KA��+Z�G/w6��B�CR���&��d�}O$�Ǧ�i(�z�@��F�V�b)�'�i�C��*�������F�j"�:�!(!f@a\�1��O�) t54R�B��B��,{nB�u���3�/�t�2�gǐچ����z�@�:��=<|�k��{�SL*C��uz�l<��d��ly���y.�Oٽ�&�GL�gm��@f��p�Z�b��&a�؉K!��JʕB�\!8|MTG��-w��w�(�`rm҂�_wk���A1hb_�WP�����'��3��O�GMt����>�@����;��*f~d�g�j���P�-�Xҩ}s�M-&��@����$̠��4L�Z>����G���[������H#2f���f/܃�r)��THuH����H��<�:pzT��[���XVRd�NIm�6�Y<E5+����s�U��f���Ay';���l��H)
&����\p%��L6o��F֩����m~sd�Ќ��F��fy�ͩ�p�����͝Hڻ�޻���m��o��p��p�t� #_�?�U����������<��PU%4�>�����R��^��Q��;���[���X>�3¿R�oV��z��F/,lV6�?�Q�S��J>[_���#�N�(����nJIn��K8��	c��b���ħƉ������/$a��/M#zOҨry+�w�a�4pf��~�7��9!)��8n����S����l�8Ӷ�n6� �\:!-mA��v�T(8��4i9�dBB��QGb�b���e�.�w��kq2�}#B�b��׊�Ȓj����q�&�GB�o�e$�Y�������S[P<�Sš��9�J�����u9�n�⦾�(����<�
e�����gb-2��l'�P�5'�p|�Nڷ���]�c+���wm��
�M�1�u�;�v#�U�ț��%���.\JԦy�݇����5�%#dy�e��F����a/���>�cnǂ���>�q*��
B�,	}3���ϱ�1M9GSegɡPH�[�U�\ew:*}�Ж��� jM~��+�ά���
���P��p�Y��&�"E@>���f���1(�Y>��6Ծ���{�>���)�e�ba]��@��D�����%J�DJ�]Ҩ�����>��4�h�M 
�dL��b�.�����Z wH����;��.٫���5�|J��J�;z�c�d�l6�7g_e��0R*�3B�+(�*Q�"��Ai"s�Z�)�g��C��S��Ak�R�x��x��l�!�U"=���w�5{�����֎%��5�V�(8� ���;�=8�6l#I�f�	�s���B�|>�2. �͍�C/3i��P֒�˹�QiX������zO�cq-�++滘�~��D�)�T�`�J�������%�C� ���,�P�9�l[I�!ې���7p���)�Ȍ�&����`8���Z����n~�� [�_�
�Em��Q��<U)��Q�R��Qr"QZ��h"�Gj��.��
��0=T���h�yB�KTow���~<�QŻ���*�ʋw,�����$�;$�]^J�P�|�s�πds�X��1��>e�(����n��h0���B&�F���煄�z�'zv�k(?H;����w܆+4B��2��	�}W9��6����5�6�8�/-�9%T(%4��B��e�����N�C�^����s�	��$�r�7���R�^CL���.t�8�-�-�\S1&U��ʑ���%��3��M�`���Y]Ht�& RtS?���4�ݽ~��ZO��\c� }�eC+��\~1GŻ� ]�a\�+:9k�v��\(�`���4��֒�d�,bZ�6t�bdK��w�	I�tFW�$=���=15�0X��]/�;�eQB���V���~.:%��k�[F;�Ѥ8�5]���߸�.lt�����t�q"%�CD�CN�>�n�t��晕�`v����������e��ZFq�qpao�j@���?P�%@�S&��Âz3��d���3�ϖ�9�0Z��+\hX�(P����[�h�!��E����6�e�;n�����r��e�� 1�Op%CO�2yT���V{J8�����v�oѮ"�Rb�V�s��_�u��R�"ǋp�C�NST��Ȃ>�n�U顋,9F�%�˨[J��_�_����w� ��ø�~��!��b�����Bh�Z��|<A�@��s���b�~8,_3=Sf,���"�N�f�S����9f�-i�w��8FS.�_�xx��ۆ�.4�	f��6Au���n\%�=��;,TW��EG�L`Iɜ#)�ՂY�����.bȈ�����X����3���`s��ȩ�H�%�����ٳ5I�j_ś�]XkQ�0(+��9FaCN�T�����rm2�
ra9$[�ѺϏ�s���q�z0~N���X��&��a���SʿxBrܴo_N9 �n�	�d��J��o4,�,�17c� ��a ��� �w�D��M�;Ƣ�b��Śk鱯/s�8$_v�`���W?� �%"�/���`8�~+~
���ڤ�Ʋ�/�'"��y3�<����r8�'.�^���k��b���ˢ�~j`��"�K����F-���Y��9DB|>m�d��|#,��sG���<�?+0���)���@V�+�.��
xKV�r����ixmt,����B)���=��/]�itM>/�ɐG�$�7��7(^^}[��{�id�.wPU+�dY���]�i$��/�2r��>A�ӐA(���*��m��tòBN=����	���_�?�E���tDS��.�u=�Z@�/�ѥ�?�g!]l�-/�� ����atx�������?RQ�ߦ�<����A��;�C6�tB@���H�[��~�,D�X�4���_82���s��r-T���*T$_OI�{u^n1_$qw+y��0Ch�O��1��Y�օH�|i(��mA6�]���mif�_���N���f�RY���f���~0{.��;0��c��{c-��
��\k4����2�j�(� ��9>p�p��G4��D[6���0��K#��D�yu���?u@��J�i��V�d�n:v,�;ϫ�������@iL \���(}���Ŕ��;φ��I�s�m⠙jfw->.>����>ϫ���٢��}�>>|�	�- �P��k�4������E�� BIӝ��pZƋ=;���2=$�{��� �ẉi��M�.��Y)9��EZf#�%P�����$Q=�bc͞���\E��G3����e�^��\�c�sF� �ܲW���T@�sK~�~^�e� 4����}���n��݈o81`+� V�_�|Iu2 �ZΈ�ͭ"yI������V"��p'��	�0{��s���].�3�j⋞��y�u~��d�?��&1�		��V���+�j��m+}a��h@P��EV�7Oi��k����村S�-L�5#:��� G�E�2�FY�fl"&���W��V$zG�����u>X�gß+���dd��-q ������ͣ��p���Ķ圜 G���'��c�R�Ԇ\�"܌z�VtLk5�iV���{چTr{���Jg��B�J��o�'�ͺ*�����g���r(��`d�kvV���B
���<��,��ZYRO ��H�ʰ�����|R��}�-[G*b�{J�p"��:tw�
���Au`�L�wз恩z:Ծ�
���'�g�X6f�<�*�q���h>=�]�;��c�弳ʩ����4������`�����W�V���m L�V�sB���p�;ܦw��5�w�mWx٘e�Mߝ��4�H+�~�l�I0���?fC�ܴ�F�S]'��#��ί�gy��D��ߨ�q�g�����Ε���$N	}� �f��X���2p駫�_��Pj���ըO�cI]�����cjm�_���(n���C��'���AǱ��=x�����S�1��k�n��u�5
�k��d��i��ýNJ�,{?�����z�8ıT� �x�!�@���X*��	�lgƏ�9�n���@2X@T&�p+2b�Z��E��E��g�+8�}#�Ȩ@g�l�{̸�<A�����ʹuf
s�t���C�-S��]�W���!`�;���@\�#2	v%J-Q>��0 i7Z�j�R����\҇ќՒ�hO�>|���<��M��c�4B��Xj��	Yu��6���%��J��?���08_`QD���9j+�a��d���
ȀN[.d��OTvљ-`��o��p2X�u8	�^N�ve@�q�i�ri�%�1�H} �hցb/�6u���Rse��p��ć��v�I�E�@1�!G:	(�7zt?�i ��c�=�+/j$	�]����ʖ��gϑ)��n�796v��$b->I4����nGi�il�4N���WU�P�)]H)GW�;���'=K�HӤ9Dc˟յ��C��>����Q뙄IK��)pꑊ3m�����U#ʑ��!҆�(=V<���W,{���1u�#�+W��#ԭ#��T���@�S�s�*`���V�5�keB��{Zԕ�rK�kH�[�*��y{e{e],���p�v�)��v�ϑz�p�����a�a�Ȧ�-�T��RL�~�����C�0��P��`���<�9nd_����-��i|	@��	������{��04��~%(���W�@�m�^5���cq�� α��HF��9�sdtN��^2]q��gN �)_K����.RX�D�%C{����S��4�h+	o`���D �c.X�>lVFM����2�N+~���ч��|J�@���fE�������+����_���Q������s���^��p�������~���{%#���^篒�/u�����OL�T�9�{a��׾}XHs�L�j<[� ��-�"Ɂ$�%�GM�Ź�mp�l%�k\�г+$�.=���sF�o�q�i�����Y��[��
�����TM�����I���6�3m"���"�c&$'	�^d��D��W�R�^R�Q��$�
$�����|>k<����9��T��4Y�E�%����֠�4���.�l�Q چ�	P-���#�����\Zq��ow`8�l� X�$���|�ب@ι��^ތ�Y�\I^=� /)��C���c� �|~����p���+�dԺ��7w�<��x����8��k�␍/�Q9��i�zf�h�U��/�N��� �Ow�o�S�-����?V���:6��S���s9�`"�
��Ȧ�?��V@�\q������rG���l ��b��u�����b����!S{V��X(ן�ѾL����b!j�9�A������0��8r�{�j�Ѥ�NB�N:�$�u�%syv��
>��� �)����JF�ϖ)�!.�:>�8�f���� �}��TwA$(���?����~�]��q�h}�$���q~�T�>A�~ڐV��L����p�UR~�����w�c9�ȭ�'T �cH<t��2����q�d�@Y��2�b�n�ÆV�ъ9d�n���gCOha�AԾ~���t��2{�n¶�F��_%�*�J�o�O��.�I�gOG�	��i!lOc����x#b��A��_TF��E3�-kz�/��}���?�yTä�~_��72F5L�����z�=�J��XD���2�N�<ړ�;�F�0@ˤ��� �&g���!X�n��OT��W�6da��η�ߑ�h��a���ŭ��q�\�ӫy�U	bw�k�Nu�a�75��ٔ�DZ��x�D -}��ҭ�d,����d�Pa���?]]� ����[C>r1��1�
����~0sh�v_������BTۑ��$��|"İ�I�N<�Y�/�o�7���l_���!�#���E\��)��������f
�D��j���!����>�<q�A���uSX�ݦ��#��c��}�xCx)C��6����ዉ�����Ą��Ro� I��t�1w���[F*����������I�`T�
�G�E�t2QXr��,�(���^�L��*��,�z��N�B���k�˒���=����a�R�7u���+���H�N]�oI��Q.��N��
��Qs|��ۛ���J��l�s��g���\�@�'Mu3�h�Ê#�77IYx��&��
�0E
���ZT;��w��?�wS���XXz�:�H�UYNkm(Y+�
��.�3"a�TOd���'�~�۝�������J�u[�1����%/��1n,�v�V�;"n�z��}B��E,)-���u��rҎK2Kd7��R��A���=�x�N��T��8�Z���Ͷ��u[L���-N-*�J�XS0�Mo�C�*�$�+|櫖Y�g�S����]���Ni�r��n������%Z��wӒ��W�/�����#pWb��|�\��������w��Я������B��f'(|u�"S DN�3tz�X�`�����w��y{�o౦�N���Pw��Q�.���*��b��u��Ch}B��$��Bx����l��0c��@9��y;n.%	�OE�>��\���ˑ��S8�AZ:Tuv��p����5��1w�
�����Ƌl�(H�b_7Ҕn������&�;�u�H�V$�E���3�ڇge�rҁ.X��b�֢`k�]u*�@��N8WZ<��Җ�͔�Þ���C�1�I�I�u�OC'���ڼ;}�&�O����ԧ6����W2���/Ɲ�KMW6՚����NCv��@�I���ox:J0�|�`ȹ,fP �E��!a~_W_z���s��,r���w!�A{0�?��G�Г�o��g��Ͽn{���Ճ.LYG㸮�/��ˀ4��rř��-)�F���_�(z-��Z,8�uƮ|�eE5�XG�ɏ�M�K��-��|N�������Ssn��Λ�����e<��0@]����{��A	|�D�J�(�R��$Y���A�Q�N[�"m���󦁓�n� �l5O��VƯ仚��C�:ּ�oM�z�d���͵�Vr���jb�輩�Ob��F��&���%��,���Zi�yC&=b-
��NҝD#f��u���ڇ���k�t�c��N�}��8�Z"��ƚ�5�y�l�C�N���E��|����ޗ����T�����?s^�=;b-����0&�b���l��W�qP���q�&fuL���0egA�)�q�;���Z?���%s]A+/������rq���-U�C�4��&��#9��8����e�(��ۚ�=9n��$q.\�$�����Y�蔃O0��z�u��ތ�:/G��A�t:��������@;��I	�a������ed��YIۥ��{z�ss���ihİ�4E@O�w�AO�\U$"����K��I��M��T������[pF�g%<��>AX'��߉��X��fQ�s�}_MFґt�/-���
��\�e�~^9�����D��Q�����^Av���c�x�g�ΛU�-g?�s�4�3i��p{��r9�cg3ҧ�%�!e� ��Ibs���@�t�����#yL�İ46WR`f����Q~!�>U�@'����J��֒�[��M_��K�����5	��ᤛI�)�Ck�p�B��Q.$����ߚ�fe�&(U�o�������S�4��k���d��;�W���^~�7wt��6�l�K��qYWWX��u���Q�y���;S7x�{��������Y���<�w%熪f��&ߘ��P"���� RL���Q_U�T{F�Q��	�IE��շ'�n�#R�Q��{B4q;x��
��N���Ţ�]�Zh1y40"ֿ6&�]�D�U%.�X{��=m��*�k���Xp�#%f"��d۾�܆d}D Q�;kCGN��H',1������S|�ъb���A�A��*�C��o��\+�d���b�7)O�qJ�Y�|$���O�c�6��T��1C�{����1@x�������M��⋘�!��{5ڣ@��{_m[m��UK�bOTX9D^�@L9�ae9
��K?�O�ʟ�2$���D��	P��ORi+u��m2o�Y4�3��ߌ��ܯ��Q�̼˩m�t�;\脐����w�q��D�����?��8F�WX��{9ac�5[�	%"X#��^Z��BQ�
�7��{������4�]s���7<��+߾%	h�O�ZS[�ݠ�{�c�y�7��ew%6?�3�#�!RR��!�A�ӆ�J�&�>E1�iy~�����g������������5	�z�Z�#��n�`��������UW���Ӧ�|Of;A����{�`��4h87� ����4��"�k�k~���f�� �_���/Ә�E�y��ws��t\�O�Df�W�pmYJ*���T�ާ���83".l��<��v1*co9w��b���^{�9z��[�-��GQr�]��!�bWo��Tɽ�3S��EjhfM�2^$k�Ҽy��|Ж���\�.�ϊ�nN^����o��Κ��a���a"�C�����Ԩ�UΆ�4�5Hl�Z�O�$�-�٧�90�Ȁ*���WXU�E��&�~������_�+d�_i����~�>�toA��Va��#���h�!��{W+Tv`A�q��ih�V��M�A4�PH���O��fb�!Ϟ��).�Po�`����'����QL�"��w��Dc��ֆ�[&�:���V��ڹ�<�/J<ٿ'7�c�'��¾&����=)���`^p4s���<�JF�#l�IY���ÒY��0�N��ݵ*k�(��f&�m��"�m&>TM��\�v`�X�U�������aE�Mȧ��K4f���=Mp�C��.�1�C�����@V����V��_b��g�P> q\Х��`W����a�]��iC1A�wp>�^g�bo�A���"�gV4'TY��7�j;a�ȑ���#�9}��Tm���=A�ϼ,F86ٚ1Ȍ�,��C��=K�2C>�c��b�0Fi����j�3_�!�4C�=U\�Ch{���'{�+E^�e�MO���hh8�^ؤ��X�<r���∅&2b�R��:/C�4����<���c���B9OZ}OI	�)�����4ϋҭ��~�L֮�s?������%�	;6��sg�?X!���s(Z�f���ܢC^�������$ZE0z��3/lF͂�'ē�-�>w)��إ�����`�?���>e6*J��|~j<�9�(�`��3�y�Tż�5	���+�
�Ӝ_˜&�O���<�
<	@�p�����i\������������i���Bb�l�[�渭xk�E?ִX�=Y���ώr��������Z�Hɷ��s���>��?\}u@U�����Cꒂ���E:%�K��A@BJ�J#���tJ#)ҩt���>���?{fwg>S{f��"�]U�d���{J��ّ��ٵ���ϕ���^�a�{č(�H��u,��c�O>�i�Y�����;g���|���5��8y�@�.^r��.���5�y�9���冟Yi*c'֤���b��^,�C
D�J����k���\���:���ƭ:]μ�73oYeR8CkN��s6d�1Wfy��_�y�:d��Sq�}>;(O��eӶ���FQ6+�z�C��Do���r�l�\�~[EJШ��#]�P���<v��-���},QԒ�������?*�W}}N�7� �L��/�k���Ifa���r=�ߐ74]�+��%'���O:SF�v���"��� kƩ!
�<�����.�S�Y��z��&�'+s���/�~b�����W&�N�y���"��&1�t[\� ��{��g	'٦��Û5��ד-�@*�1��px�h5�Yޤ�ў���z+���$s*baR��|�B��<�Y&7.��E��y��WK��_�_��	+��������*���̹"U��m��)%�.y�7�.T��� [��|��@������J��+0�c�>�t�J2&rȳ�K���`mN�O��ҋ�<w��v��\_���J�
Pv����N�t8CZU��J�a����-�L������r:��#�, �˖ok��d t�����VdfSғ�*<f>���?c�"�rC��������{�[�%6��Zh��X��°�2��:�!�喯Z�(��+I�}> S�)k�.2s��L�c�1��ę	R�7���__J&o`&���o��+k�K��r��t&<|Z�����$v��GD���k��qf
:����^8}�U��m��jS���^�f�[@�� , zϙ6��Y�h������ֵ� ��H˖{������-ky)��,|���e^�|�Z_�%��ن}��o�	�XT����{�¨i�b�m�����q���\s?�ٱ�~K��*��1����q��x�Gd"FY�`����	�`��BT�]=F��7�'3����b�p!��b}G��];��m�B޻|/_�˰g�uq�!&%��wC�H���4�oVx�8���tnؐ�yx��y�5,���Y��M�z��Y���0S��T�b�������F?>A�u%���h^���nm~�v����R3���d���{�jp������� �,cQĪ��n��O1�.�E�#����~�6�}wfF����.1�;g&���y<���?����fSج����/V1�U:���.��G:X>������>�^oI���Mx{"�˾���Љ���=u�a�n}�(tALI��!|�w�s��<h�t|�;l]x���ru��<�f$�����ކ넋ll���z�J\�=�T�.����*�J��K�%U���fz��d��~�X�y��u-��g˅�kz�d}�ϭ6���w�s��T>]Rݬ�Ni_yH{������ɿOp=��G�Q�t��ryG[d\�n��>Kyu��,��)r��wl�n\p���J�fi�ތ��XՖ�-r�Đ��`L ���! AeߤБP��l��7��Lfi|�)AX��-Ҷ�g�L�8�ӣ|,�?/C3����Fp�O#P��H�ʢ��}eB���^ � L�L�� ��l��N	��5Nr���=��m"��s�Y7 >�\d�?ʶl�<ߩ�f��֩W3�	���]7�N֦u��&��@�(�Q���;�.�vV3~+���Z�i+� ��5��O��ܘf��bKXr:HI��BY��t����4z���T����˦'i�8�|�
�37aX����羬�R�7�a�}/H'��s�����О�J*�|����該��=�*��/l���I|O��ZQ|�L�ʅ�+��-�~Sv�Q�&g��H��)�}�sr?k�A<"�[��RBZk���>�N[�/	6">�X��Y�+$Z*�WJ*�T(��C�Ƽ���I������՞VgVm�/_��;����7��լ��g�����}�	���:�V��p�%䢟��K���_��'ۛn�bMJ���e]^b*��6�!��'	5\p��3|,-��dZA�S�GWp}�~���U�G�O%�2�����dd�bS�s\!bqqKq�:���m|��T����������-�,�_!�8v�\d��w�d�p��ҀO���D>w��5��
*6�c��օ7�>b#�����.����]n��[�V�m���!u_�`�.�%��#v�u����{��%�����54D!��DF�ؼ������ٝ��Q[�g���RRZs1���f�"��?=�F��VOP~�K8B�\�򎂪FR�ng�^!hSt.^&�p���~�����������Z�t��U7�*v���̾�f#�-����y�u6 �0]�n���K1q�����S���*����N��@>����HK~�������3��mpK���җa?K7��8��_����=�m�k_�A�2������X8��.�)|Wh��*r[�s@N.��V������.�hx��7=��k��G�1�D<V�y,?�f�b7���e���΄1�kv��ջ~�$�興:�P���R!��<�&��A�9Ӻ{�uZ�Vo}�"�;G	�NE��d�Xpy�5��o:�R�	x�wib*�Vp�d���na�V�(�.��j�O�L=d�qpR{��_�E�����*��˨< \��
Eq� �RBW�6��v�2r49E'n��}^/3(��CW���N8���T���#��l�0捍��	�ʬU�6�6��T���zE��fI��kA�sB06�rcB<��I��[���1�;�E���ḍcX�¶	4�8�~��RWy�4�}fJ�ź9��ơ��ݨZC>�h6�Yޟ��Z\?V�}��SǞ����\��~��" ������|��k�:���Ͼ�����w�=k�J�}^�4�NΕ��ϵ��g4�rwRJ�k݈[F۷:�<�WLR!-+X���Ǽzb��	�R}�u�/�9v�{�M	!J��ɦ�{�M�Y&Ɣ�b;A.a2�f�YTe�3сP�_Q�����h�����������=��e�ğp�B���6����L������Ul�3(fB �r�����I�jB�`i��f��C_k�d�^6��ui�=�h�ρ��Ѐ^�-�=��D0wNC!8�`R�bC�I*��� F�Iit�W0O��T���sW��+��'���m"h2ڼ�^o��l����D]�ÈMMpc�1�WDLe��7잌�8�tmF4xZ޴x��i��'��� ��Y-�!�\�^��!��D}�㙹����t�ݧ,e�5��A�=���xl� �R�{�$o��{V�q�,zt*o���7���ڔ�����ªz=�'6E>pDQ�1dS�����s�]N�׺��z!����L`��
�f����4-�)��sO��X5���X�t�VppЈ��7>��U���V��9I������sz�B���B�DS�r`+vm��"OmE����D�2#{hZ���k����TK�	������+Q����H�����x��􏮺/��j;�?�ʘ�b����U7�0W����&J������ZP'����=(������4>>-ٲ..�̘�0�M�&�%�c5F	K������c�̟�tӘ�E{Q³��	_�BS�y<锦��#��5���GgZ�|\��:��Ѻ9%� ���B���h�1���v���*�I��?�i��7y�N.�A����/؞zv<�)�<3a�f!n��syM6�͞�FK	�I�_rS�'N&�1�a0��OI�9��Ӆ����ヺjĿP��� �G�����|��]�)"�)Ȍ�E[���]�	_J�&H�\��D[?D��TA~�[F96���}��"M$��(n�dNqx�Q�i����+qK��W��h�܃��c�Vԍ[$�A��0�z3?p�\?�Zk�v5(�0%��6���U:i����&e�#� y�Ρ��D'WF��fI�!eb�����(����++�W+�ѼQ�������D���֓���p�cx�y65l w��Rk��f�L����]���?�M��K�E `5s%Ϗ��x+���E�&���~7�}Z�E���A���Fl_^�.V��8�)�^��Gɧ����W��&J�-YcL)A��=>�=b�������λ�K���oR�c�M46c�8�+!'�N���N��r����0Q�BS&���v_kF�E�;HBIFS�a�^���n���/��4���H��	qs]h�h���o�]����d@t������_�6N���C�G\���#i��H�Ӆ��,o����ʠ�E�t���G��Ե���� Q��Ս���� �N�ۍ�˦��qm���V$?��:�:gAE��6x�
?��}�7���ړHD�t��a��)�Ay�5�ݻPlp�����.�N�)0�|�2��y�%�i(��� 'ʕ��]y<F�2y:��j��Siʇkw�ǌ��a��Mw]Q>��$E-L�A�-CK��ZN&��$e��?G~~F!r�q�^�T�-~���̎�?07�`@�O,�L;H�6���:{�	�O�F�]Q2dV>��`�:����JWM�7S��*�U�N���`�{�?dG�ąl��b8t�ʭ`�)�tvZY��&�£]�S{/����U=�y�-�j}�׽���3A*�BN~9�)?w��ـ42���"9���.�8.n��ۖ^ XI3�\$���T��LΙ��*L��()v���r \�+�II��?��<�����;�-֠����pb֚��%6� ��CV#� �~�%f���X�b�{�����[������agp���D%�']�$x������K upϦ@Cv���u���h�:(���#�y�'7�|�XOZn�T����-��A�3�t��U�6۳��#Hp�o�&��(|�@��ӆ>sů��� �^�yZmJ�����k�$� Q�zt�g�:Q���=�_�pĦH��h^Bj�쪢J S�����{eb����S�i���*����i$x��Ł�Mz��k�cL����b���U���sj8����t*���%�`�>[�QOxĎohkK��3ڡ��yD���=bv1LF1���W�O9û�n"0.	�z)�c�U�u��v�-ı�����#~�BC�֛��7q�p�KRgt����-���G<-~WG��-:�oh��e�|��u�*{M"��qI��~V�3ad�iNDH�ɞd�Q�]}@�)a0��UI:q�;��9\�!5v��� �ֽ!ܕht`�388]�%�ʶ��@\|��e������(��!�����5H������X0�ڂ�%d�g��BvKt��|w���'�7YV7&Q���o�u{�I��Қ�@�!\;�B�Wkn54���ar���L^5=�t������C�l�9_CE�O��-1�ѪK��K�ڱ�T��n�]�z3�����*�~����v���PrE��e#�2�5.}R�Mm-���}_AaZ���.Y��������Y�Ve��SD��X�qQ�#���P�ј"~�?>F���^ #r�z��9�e��I0kYb'�:�7�)�dsE�w7&Į�,kp���s2��T��ŗ��'6ş��cU~.�"��I�S�b�**SB��G�Lt$H�;]���B�
Bˉ��v�>�r������R�iMB����۷ 	ׯ�2��t�F *"�I�!ܺ<�K� �"V� |
2�$��� �w�p��%�R���CMv�����J"jE�b�ď�?G1'�B�G{�0�G��#���*K��"�?���?T��6�?�M8�UH/~��59���57��Or?k��3>O6L���D���M�D�(u�(��:��fr�K:�!��V��8��R�G�]+,��i��5�3&�0Pp���<:u�1���+ }��|~y�� �j>kx�ӛ������U0���ЊɄ��&���al\�4ݰ��CƁlY�0K�����췳U��~��
���X�s�*0K�?��0�v��/M�d8��p�9�l��cjj��;��'H��ɾR#�Bh<,n�ҙ91y���s�U"���Z����GD��r��2��c�vSW���)�ΊD��:{�}c�R��F�����?�K�+�(rb�N!��a������3:[�LӾ^Ub���2訖=Qq�s�_���ya�k�N�i�/�<�?FQ�џX�N���
i�^�co����nyGA\�+#�C��K�F�7���gl�dA���cTAl�n��~5�BzB��6�"����1���ZJ�Q�V����L/�,T��ߤ_?�-�O�
�{��c�i*�\��Prv[EB�a{�ߚ!Pۭbq~�\q���w�B%�����8�A���fh��Vט��RF��Y��H��f�;�)"0f���栢������p��2�P�$�?7���C�o`@���&�B6]�<@Kc�xfI�x?�ц}}1�9U,	�$�<�u���u:>-.�L��ᣞ��|M:��1n8ls�b�<��-��R|����x����%�Jan��
�%Ww6��}�ѕ'��9���+Y�q~�:1'7���y�CH�.�`"�\�1��&`Ȩǣ*Ӻ����9���ݨ9Z�z�Q7@$�F�x����w҃��y��#��Q-�m�u~{��A�r�P�����%R��O@uafU{x|�q�5,�wqG��2l(����{/�	W^p����0l���}�Ml���e���9�5�0���X����t��]-�#z�4z�mw�L`;"w�לY[��Y� �;ZZ:%��J3[%	�����6ƕȊs�g.ފ��R;9/]t'���6�b����k�W�)�%A�}9n̃o�?P|Bi�Ơ������V�bT�-�c��WW��*����6t��3�o��IԨ��,3	嵝v�9�Y�^�^T�5�%;��Z��:��cR+p��YC2��)"R�%0�+>d�Lڥ*N&�H���
�؋�F�o��H�j+��<��7�i�͇�Ryq��,�T5������P��nIF	�_�!T�*�(U��n_,�ۥ�F�Pn(mC� �v���w�f�m�U�1��柋a�֩`�i7Ó�w^�}��=�a�i4��N/����k����!.=O`:HS����dE���m���F�0�&�Z=^w��y�����/rZ��(�7Z�M��=��Q�!ܟ��F�#�;<����gL���d�*�"�z#�g���)��E�^��|z��^�^�b��Q^̱P.�����J�ʋ���}ܻ�8��}�8��Ti�iG.����9<���Fpli����3X?���FY�aB:�����rz���!��lq��C�*e�f����e��Z�^�Xϴx11:�"$Sz�'� n��>O�*Hd��2l���<�q�<Ú+0G1RT{�-㋶z��EW-{������/Ԯ��.���blA�q{�K���S�$Ƀ�ϫu�  و�[m�io��\���Ĵ$��9��Mւ�`�$��XzM�mu���*����P�j�Y�aeBXX��b���yx�z�%%jY.���r��c�?�#�]�����-B �%�E�՗�T�<��Jxgk�
�M�L����SU�jܾ�Z� �������"�������9��4GSB7ߜA;��9�eͨ�BW˛��W92K��O��F�<���Y���cz|��?�$���Î�ý���c�]�(��i�A���}¢/a;9?藨հK��f.׸%j���3�}�F��~�� �<K�8%�B��'�7A�>��Ԥ��;��St\0wC.W��#��K�W�E��zއ�8��REq.��A�c�	���-��L<��xJ6H��]ۮU3TML�V{ź����3��f��K�0�ĔG���'���[.lR _L `���9��\�j�I��(����ӭ4)t���$q�@�a�	� ���n&��Њ~D�V��ݼ�v��e���^�e5~ݳ�~=�#t�	A�]�=	3���Cq�ى�w��7�ʻz�xD{�	��WG���nF�)F���G�L�7��\E]�p�,wG~����WL�g���ೋh"tI���N|��k���Cn��a15�P�2߰ Lτ����)�s���¼vߤ	�f7�7��+��1Y�Z˾V��𲲔���_����E��gS��P�7�l$(�Qq�|�O����� �����j`cљ�'+LO
�0�����i�8�h�sٽZ���S������|�:˧�A	��Db��hy㮅��rݗ��aj=�?�ԙ/��+IA����'6T7 i��qO�6{-�>�R�~7)�0���0��o,1��B�������\�!���#Xb��P���?Z�m���>�r��a�D?�B��x���I[1���3V�I̱�����L�&CW����8&B pW$P�r����&l�����1�)\����ѽ#!r��)�A�i�L4f���S<�MV��>ۆ}ht�V��U��	��!��zy���kS�nt�j{廰����i��a�RD[4� �'�kh�	{��Ź�/�!ʢ�<�5^��D.���@�Q��o�r��w9,�k2�\<�=�/�vIΡ�8��9��%*�������v�o�[���w�]��s��=�a_�N�G��2 ������9��.��f��S��紦��os*�>[L/�߸#��.���� ɠwݪ�A�h�g4�( ��G��
�9���I�A=�� ���\,��޲ �PV�|��D��d�_����|B�{]ks�ԟ�݄�L'�O��4�8���G�0F��zs�1��J�5"�!����҂<�_�>O+5[ǘ���{;��-�0��-"t��VDƈ��V�8,�vT��y�Df���-��z�M���K�/��k�@_����+~�|� ��[\�M��K��#F���c����j͹��1X�q_�k<�<R���%��(�&�����6�]��<+�*e�<eok�w�;��߼�Z&�H�ؤ������nW�o��KW��ܿ�j��Ĩ���@�J�i7��	簃+J�eל+�4��2��<�,�6�PYqb�1��P���	�pkB��ư��Ⱥ	k
v![���������	��NB�ѐ�ׂ�Qx�_ y�e�?H,��[s- �+l]Fc�q���/��s��(q����"��3��Q�/[t��Js��O��o~�>;�*�#}��pn�s������`�r�1܍��~	�S�������V���dO~Ò� )g�v�<��wm�[}Qv����=�E���-(��?�Ru�Xˋs~[:)u4��K"���2C�F��\��s�~��/�����	���A4��3?����8�Kwx���YN/�kl�i4Y��^p��;ia�ϥ_ �	�jҠ�G9�S�+��$e��!��۵1�h����W�C�/�&/L�͖�ʉf���q��{J0>DO�\�!+�% M����jZe���0g�`O�41��ym�T*x�kL��^��GL�s_Ȟ�������0D���^x��xk��g��#�Ñ���}cI��YN^�o2yn�E@�"K���������MM��-Od�C�A� "d�|W}�����-�W*�Q�r�� �<��.��]���Q�3�T�]au�zu��1�?s�x��0Ϳ��Lcb2X��)�gX�U�0s ~13R4�1�s��+ZĦm�e9���,�/�}��=mN<���#l*ڼI�,+�M�ٔ�h�4��g,Ѥ�5��}�y�G�i�qO���b�,���h���]r��. Sj�s3p�p/�Н�-۾{����m��7�8^������t,�oZ�e��kYP���R&6���n��9S�"��02
L�N�����kOi�e��J�U?Ȧ)��<��(
$)]�`��1D{Y,���pN�r�&lO��� �@(Ya�S'�*��1-�����|]@����=n6�riK�Ș�ڬvi+�D�m�҇�q)��&#�jvq�M�!�CN+�)bP+eN��fR���=��c�
<Ǚ����*���Grw��7��D�ќ�ww�z�P�пy!�{ӸM����*5TwH�*��iZ�#w;k�6}~'Ih�쏀�<r@NRfD�<;;!�_����?7�j�c�7����F��yۓ��/+xT�c�o�j����kZֆ�J
�k�_q��l�v=��G��͘m8`��������c�+��f7f��V=�˭E��FT�.��k��څ0�w��,����ߦ)������['�?�RV$��C��y�E�hR��h�8�$�m$�޳��a��1d�z�E�;�9j����D��H \U��m�{���v�G�����I��H";� �H�u&#7�v;�`g�ny�?��$��}��2:M�!������-�x0��HD��*/k�2�2������߻���F�h���M��
tJ0n$�W���B��w���D2�o��ҮF��?����Գ}\�\��^�8����QQ��;!��es��;��24b��XY��9�ϟ�9U';��� 8(�O���>���!��-�+:�m;a�W���\�$������oDRRgm=7:�]� ��*+a^5�Ad���IV�	�D�Jpt,��K(mԞM�^�ɂ�����}�(g��bnL3��g.��7�
������t�y�����CaV.T A�o䒼��T�a�~��:�Dl��%�Ǵ~�w�éc����C���x'�"�]�{m��f""O�
d]#�5\
�8��5�\\�+%=�y�m�fՇ[�[d����^2�X�tzr��S�w^�c�	����d,Ee>�lb���@?�|iD���>������W�O�E�b��-�yVA����}IJ��[��mz�����u=�WWNc���󵑔<�ئ�왧�Cz�A������zgU.,v�V�D���'�#�f��	E��h!5	ހ丩���C��XB����hd4�J?�����a�;'R�%iφJ���zB��-C3�M�p�����1X�9�e!H��v1���8��q����|Ko,�4����6ػ�����e�H��m �'��17�nCA\<�ҧ�����5~^3O��s]t�].��
nn�n��}U`IL�6=C?a�ᅘNLG�E��d0d`kDl�WE?��@�@�JO#꽵�ϱb`�~�M	�Pχ&�{�x��I��V
>�;GVn/�FD	LˠV^�v�q*"�߬P��R_8#٥\wiX�:;K�9=)����z���B�C��c�C���D�P~maΧ�Uy�_� ��K��Q8�j�r�����wB�,������X>�N�]�MLZ}�< �<�P����
J�>I��B�t�&[��%3����V��Nqѽ/��y2[���K���%��H��w[�'ٮ�H'W�jh����ﾼ����SUCcP�����m�W��hׅj��_�� q/�l=\�^�[�O��9!�{V�<=}���x9�Y&���p�>ۣ[�/2Fk֢^E�Э����Ah��Y@�L�O�e�t=�;��*����~\�$��C�y����Vxfc=U 5�~�� ���E;K��^������~�|ǧB��V����&�|�N����qτ�<w�̻���oj ?[o��T��X�=�G�ظ�S4��}6t����yL*j��a�OHl��|#8}��J����a#���#�lW��TK@��	*�f_�y��`����!ˋ"�h���r��Y��-��;$L�|g�>�f�t��q��Y.��ќe��5}�%�N�� -_�h�u!^��ׂ)˭��I>Y�7<�c}��|b�$!�8�(�*U��y�d�U,t��(ܣy1�q��9`�G��r�;s�����6��f���^�,a֐��k>�s'5)�n����\�]Dޟ!!ҩ����$�|���O0=��)[2��H�g	�����<t���@�Q�"*΀S!Ԥ�3�o�.�;W�F��#T�ue>AZ3%lW}�,K��t藦=���_��881ҡ�G;~D5q� ���?�職���Dy���Sk����Ib-�K45�d՟��_31i�?�;O<"�m����6a�Ju��e ���3Q��@`ɾ�}��M^��f�/�iw/2~����%��͌3��z���>vj�H�ʜcVw�g�S	�vu���V�&*q�����?J�K��CVbS3�Z�D�a�,#N�tj� �n{m9��g��������*��E��dr��y^��L���kWt���A0�/�G������m2�~��U����6*	\���&�#�7F3PB���L7G��O���q�~z0���S��>0������.5� �<|ztA?�Y��o	Ջ.��ݯ�䟤�5�\/�����ݿ��o�!�����=��_:W���վ�*�'��躿BT��j�k�'v�����kɲH���wF��y�$b��	%��ӄϕ�m.��h�������X ��Ϣ�Urg�0��w���L�g����g�P1�ޭM))�����y���m#���)�8w��ݳ��'}#fx/Sz�{�jba�BP�a5`K�2� �ˉ�\]�oa�C?:4��dYp�{�F�A��z��� *�c��}R�3l��u����"����Og���޹�{�*-K��~��^��3T�A%����Q]�7��2#���|�1\ؑ���O�u���&MK��1C̥]/Gp��Vio����zy�6Ņ���b�!�ý=Z���Q������=��N��%��"&^��X��w,)9��uF�R�T��C>��,|ks|�$e��Fw�CC$!i����ы��1;���f�ŧ_�����^����`'�����X.;��mh���TU���f�S��)���+�ǚqٓI���6|�Mk�)tGбx^��CP�#�nTҽu���'��&��4v�v�N�v��Ad�!��ax�ad�ad������D�m���*�A�/�נz)J�'�'��sf"��$�m���a@@<Jd�I���݋���^�P�}�ܳ�?�����/:m�;w	�m	;?��!���=Z�2JT�k�L_��K��;j��St�Y������mtL�fz�h��8I��N����OM����2�M�)��"���'���vH9�d�y+�7	��c_�G6q���.���3���fa$�7�Q�M�-���SZ��Ew�����jO�x�$Nb=(���?��,����ZΩ�'˂O"<�Y5�*cC(��mf�:�f�z9�Eve��L�W%����_�M&�6�U�fX�E��ms���k�[^�z(���u3��.��~��.�ɨ�!��������r�M+,V��7����O�#���o�CQo�z&4D��?y�t���b7\	���c��;�ja]c�T% !9
�eG*���`#o���W�{/��f�4�lm�*��-��������2D���*��]��y �g�a��R�b��Oc�|�_&�^K������ �KF$�iF}�јA�����Un#��u�"�&��ήV��'�O#a��'I��k��
�ۼR�c(E}�9�[n�~��m��ӺL5�,��+� P,�M���`����H�R�07>�8��x��Ѹ�� ��,̗B��oo�M|���j eiK𡹃���	�_u���[�u�>م}���I�[6��n��|��A�R��*2~�����?l����s��O��!��>�o�+uh�"�(�@S�Q�ͅ��ᓺ�K�1�#���������QB�$�J�����W��o�7�����no6���{����}���{�5h����d��4k�x�u����Hh��Px�id,(�i��?�i;)��9��A\v)����,7\*���S���<����)�9�����zv����[�5¸�ƮgɕG1�([��)W�^�"D1�%<�&����_��|B�Tu-���zBx���������T,8���V���C���,�8|w�TdL�D�5"�$��Z�*�B�z�&���.�w�Y��9#O(Aq�'�qf�e]�;���W�]:�	��?��#��_b��1Sʨ�Js�"�N��b����
aW����t��tw���r�'2��3_���=�ye�M�&����Q,C
=kyR�]|�u���ݢ�j�����<B�ǡ����lVua������5Y;<�EPC��πn��A��?��.nk��P_�a*�!��R?����
���0\cŷ��Y�5/lj�j�;�P�@���/���Z��&d����pꮟ����?}~KT��C�_}�w��lƝ�gV�J�h�{��r��نP1��p�Gq���/�V#%`$�`��겔���ߴ��*�ɻF�d�󳍍���u�2082��?\�"-S/�j�չ�+�t�ޥo�4\������j�w���
O�������
d,"�D*���3�2Ǟh���P�c��H��hڦ�ӈ�����!���v/�v�B߳r�(_��!�'���N��!����҂����i]V���ݛ��؈��Ki��>!�� ����J`��F��n�7�@��R]N�6]��a`1���BV"�T���U7���(QϽ\�e+� ��ِ�ֲ#��~�C�?���?�[�=���a��%")��1(qz�.��x	1zny�?o��}V+��K\M>k�h+V�I����pwW御�4���Ӣ�;1�
R�F�.X�vj����8�Y����㓄�b����������F�0��<�'��_+�Nw��K�oh�i�]~���;;��P;Y�n(^�9V�h��(�g���n^��~\��T}����7��wд�k�m�(��E\g��y��ܴvU�WI����/�<�<W����/�	��ӣ�����T�Ry8g0�G�'4ӟ���PQ�"~�+�OUz��hsC��� AU�/u�ڸu����F�*��������gO���o��C֜8|�*���T#~,(*�2u麇���8I�	0ή�*܈~]���dxg�(�TV��Gl���� ���u��fJ����@h������M���*Ù\<��A'�T����$/]Y�`�]*4��['�j�2:�>�z��ujp_����tf�gJ�p�3�������o�$��r4�ɨ a)���R���k�U���4�wު>��"n��-�~	V��S�5�{9�m�S��~n�����(����ȠqaIl�i!x�A|��>��Rpk'�� ��b��y�KI�Ͱ;�^�ji�g�9��}C�1?�IS����+�60@�ʖ:�(����rx1zӾ!�^(�w��ΧԸ��b��S@�pr����)�t�� K������3�Ԭz;o�OI'�{�3���妍�
�ӓ8CK��3�u>cʔ�s7:W��.ۯ4g)���%b�N6k��K��{N�������d~E��{��Ln:=%d��8[1=
K�ME����;	�_�Ǹh�ե��OP���'��A���ꦲ���4И��ث�O�>�a��0y_�d���0�e��9���!��}!�ST�/f�RU ��X�'�ͧ{J��/AG*�~�ŕ��!̲ٴ�L��V.,�N����`���� ���P���X��x�N�A�M�J���'��i_��}%��C���D��{Q���d��K��/Z���%؟�M��yex��5���.a��߲�~��$��6
������.��KS�G^��W�?�K�>�~���=��ۑ��a,�r����~2{���	_X�0�P��NA����	�1��8�O�g�4�_p�zJ��Ǔ�������Ԭ\��i?�bZ��S���K\E��U�n�L�擈�����x��=�H�M��\m�~���@~`��Õ�g�i�_�"�V�L�����r��m�����=)v�����H�q;Ӭ	�~
>�=A��57Τ����:�'o�1HU�-< Z%��z���%۾�Й�- BX�QY�їP/�K%�gj���O �I�`���g9�` R�x��A��"�L��{�	M��0��Tx����s΄=.Q�T+�f��P������F��w��ĶRZ��n>
Ǜ�G$<%�
��U?J����bT����(�isM��o��~��}���*��4L&� ��)f��#$/�]�H�s�}1���ӓ��y�9�x��6y�_5{D��'c�!�;�mb����nɖ����`��M���rM�]L�����<(Ȁ��1���������~����K�b��M��V��)���L�ȔDI�xG,+��8��>�N��4:���^I�Zo�G���T�Q\[p�5Ӟ|��>�����<)H�1h�?��t�P���^�V�)>>38�/�<���WV�z��"�V���ͫ�E�*y�xʀ3`?\��r�	?�#���ؘ�|�&�ql�0_��ȳ�)�͐3�=��\=�����f������'�5r�8�p*e��&���WM&3���n4�ƥ��=��EU]���:���i�3�Iy� �Z��7F�gH�	؏+��2�̾cbl�e?�%�hu�6���rA���6�5��."ؠ�/n�\���ٳ����y���ޏ~�e��m�f8^�����%W�uTI�
�2��|��d�W�7���Q#�B����W�vӉ����9��--�)�։ w�٦ݥ|�����&��S��*
�<r��4���,ɣ�+`J�7�	L�"��>�^�����r>ǵ.[�X���Ѝ�D��XJ��k4�Mo���˓��C�G��� ���վs���>맜��Ǎ��x�ݞ�gyx�G�<�;�k�>$fؗ���-�	>��G�������c��Qн��x�hx�n���z�[���祵?}4st"Gi^ƿ����>�Ęn�!<*�i���ѱ4�D����G]�EIJ�7�-���k�`��^�U�K#�t�
J�4J� (�݈ HHI(")��]C�
�%�3�0���=#���_n}����ٱ�Z�X�\/lY(��7�O�|�FZA.;�w��$��e�QwV�"�� ڑ����F'hL��u�TWU�{�s�+��qG-����t�g/AަJ�	�T|O��g:���Ay�,)�(�����ܿ���
HF୽��_E��p���R�j���O_R�OT���g��>���1g���ݜ�9�\�I�� �e�������-P5�!����s���R1�c{&�r2:M*�������2��h�����C~�?��&Z7��E�m��)��>>	OoU7���Fg��*U�/|���yn?	r���G ���c���/�Xј��zU�Ϭ�2��a]Ef��F^@��W��is�W��Miz�s+��lB�.����cSF�z%=n���CR�An�����[��nug����]X��F��dy�F3|����1�.B���1j�������nW�%Ⱦ�iZ�9�y��>�^_A���[������דe��V]H��X�t|��ZE��Kq�dp������iⅦ�,�)�!S�U��@�5��8�F�CT�m�r��,���,��?�b�gb�ˎ�.)D݃�l�_O�Y	��%WO�1�\��BD������f֊�Ņ�/�e���Ҵf +��O�4����k~�:D����Cʫ����W)�\*EU��\��D�j�&|�]���KMy�͔��m�{�1*��˗�e$��;]�qmU�alg3Uݱ��,~A��5�vp�����Q�e+_#�pc,�/Z5������5J}[M�<��y��x�OF��\6U(�:����E.�')VV{�K������M�S ��iva���!�o"G��@��YF��O\o��������nq!���P̐ʕ.��\4+ox-��(B�~;��˄�}` \U[����k�TEI��y��ˀ|������77�#pdJ'�Dͤx���K��ROFCYdFy��!c�I����\�PI�:A,bqٌ�ht]eM�'ϭq]I��٩\�q�Gj;\�՞��Jѻ�=?�"��+�����v�"���~yC���U G��=dK��.2�����1B��~D��{�U���'����,#!3�Ճ*�����rt�\Ԇ`ݻ� Zm#�@R�
�0[�_�?��J�.��Qj��e����A�:9(��db��]�u�<�-}iyp����&6�?b��YM�: +��G���wD/b�r�Ju�s~sͷ
�'�2oq���L�5��e��L}��F���8d������q?����.�#�����6�������Mu۹���_�>�f;��h} '5�y�*��*����������H��_������n��
����lw�w��7��	3��6��i}��k�2O�3e�u���N�����:����"m�vI ��Nu�7����w�s�L���)��C�V�PB��[^yr)˗X��zO�&Ȍ,��U,����p�z=��չ��NÞp�rd�i`-S9����^Ď���r�aVS�!s5��4�����,~����i��wK�eR`� ]���\��ت�^y�L�E�õ������ �z=-�z\��aP��iH�� �\�U�1���ׂ������S��S&��531��ĕ9���ޟ������z"�2���Mv���U��G���Ow�~U�Bۑ���4K��D�/|�hj�]������g���a�����/���a�}{�O[OI��g-��s{T���g�nʴ�y�Z��^�&:��ͱ�Q���+c���[z=!mw�𛿱1�-����T���&+�,"F�t�3���Z2odo4�j��F��ӄ�XxD�����p��͂�i�Wp��W��� �F6^)����c��w���	��$@��}�1(3��7Yf@m��trr��ڲO�+�/��ZrOW��H�r��?][��j��+;�q�y����g�E/saG����/��_L}�Q�Cit��c���S��T�����`!�4ѽ��}�l-���u�Y�pB���]8=��>|��a��ͥ����}��gH��1A�W��A,vֆGG ��<˞��l��6���т.�+��yջ���w�[� h�/�U����⫧sn�N�M�ʛ6R�ͻ93���߮H��z��_̿�2Jس]��`��s<d�sW��3������9Y��ֹ�M9�����L�ҋ�x��� �C���γ��]�����I���9��R���j�@ʗ�Fgǃ�J
33}��s�z
�����k��8�z?g777L�455O�p�3���"��I��)E���k��F���F�L !�`��@/�L��WUUV8�z���8�C�����#� ������$�Ȅ�@Y8�7�k�$��dS��p��[ �}���L��:�U@���%�� \�OL���Y-E�����\�ę�,��:�� H����7jr}�@�]��ۇ��>��!���&��f?]3.@+m�n-3�,���-�4\�[���B���&U�Lc`��"A��h'��JS�SE=�y��'A�:�T�?������~������s�X���>����Ʈg[�E48�Z��`���ÍWq��H��W�����`���x��V˕J�}�N�9�Mo�	��%Gx��)�ռ��(��3+`O��Ҫ���]M�Ϣ~��Z}�y�<&p5������/fT�0��ߣ�|��99�z\N����X�X�u�I�gx��2���_����z���]��8��<<c�*_��5���թ�`,�� ��~B��Y i+��[�b����@������}!�S�0=��h��D�)�0���׎��A�3|��SԵE~�<��_K<^�D^��`�����C��
���$;�fϚµ����}ĽN���K�.��g�$���6��V���q���s���t0�W��Q��g^�4�&��a���r���3��i��ڴ|�1��x"�64^X���m��ϐ&>`�j�=��x����jLC�WCz��Q�D�v1�-���ũ�kG���wvvN�:� � CZ ���fE�X��|#�3��X<�k[=�����k�ͧ_�D\�����?O��x8/�JN��0�N~�;�ڝ��[��ɣ��Eq��)-������8f��<@p�| H\QQ�@J`����@�l@�>	-o�� 1�i�H{��4�X�;��UYt��x퇀Q�K�9(6��������q�����;H�L��*�Xz��LMna!WsK��yFX�<6?L���E�����2I��T�!�@�y`d
T��:ո��kl��p)dɥ��M{/��f��[Vѓ��Ǆ�����jhX틭��~���y�~�+�T_,5/>V
3p�Ó�����rw3�z���m~Y"k��֝gg?��{A�k���wW'QF��!���W�+ͻ��Nm���ߺ'Ҍ~��)#Ԅ�52��~0��R����Ih{��X������x:�ڲt媤$�:�����PB�x+��KN��
Rͫl�.V2�GL���|´�9w�YA�m��@ʭ�D�����a�?\�[�2���?o$�5��l�>�)0n3��h?���:��.��o�(m��hw�)��P�G	@��~��^f/K&��8oc�b��=��V6F^� A��^���1 
@�[�/�uD��|���G&���g��K==����� oaa`�oS���8�Rt��?HO����3s�Jmߤ�`a&`ΐ159���mx����lfB�fMol���f�L�3��:�����:##��j��L3�O�3��TJ��G q��1eg�6��(�����t�K)���{8&Wmm�_/@�;D
��J{9��dq���ބ�[������v����?a�8n�qo+u�M��T�Bn�y ��o������un.Մ�5..�S-�jF=$止[|ǔKݻ�7:�i�5�@����Mc������������7H�O+�*��Y��ζn��:;O4�&�$�P弘PŢ�H^e5y.��(����g��s�,O�&m�pn�5�,.���s�3n���J�%[��R�2���kz~�شl�8��Ē��h֦�v��Cֺ���~�Z���KRc���N��Q�0�u�������v�U��^H�e-n�	�oxJ���^sm��rrTd����M�g���6Y�W��!��5c�����H:
8�q�b̈�3�1�<i�_�mEf[�-n�O����ɹ��f��� غ���y�
�A�*�����Z���H8�R�҆4`�3�v+!�8�M�|9���,�"P�W�Ld�ᒕk�\�10hZ21�r�X�)��/rq
|����h˰ޯ�´B�m/�����"�)���.�KY�;���G,#�N��V}wd�
����~ʂȝW�_�FX��G9ۿ{�I�RGD�Q�A���X_�r�$�̥ԫlJY����|�r|p�Q?�hU��u��C�i\򳑫��*�L�!?h�U\�O���m,,sm��q���J��E����ҾK��Its�#����lW/��1�8�������?P�y���M�2]-��s�nӬ7���>�̽W�gNa�/O9���m]ʠ����������%ޤ��z�;� �ޅ��Y��v�+�G�I[
<�b19(ʴ�nwC�m�R�c�'C�;D#���3J��B�cY|��o�ʋS��f��ϛ������3y-�OieE>��L$�юz~�{aO�*h^���-�r8�+K��0g\g�|A ��/�� ��K7�� � �>���mh�b���� ����x.��E#�k�>CR��t0ا��Sʮ�`F'q�-��?El��R[�>��]�*��΍~�d�[�	C��x"B>���,�����6��H
GI�5���O��}*~���<�q���#�[�,9q�r�K�nd|������@�����K]?l%���R�Z�*'�*�^f=�����5���)Y^����?�\k��߷��T9��q���P�:O߂��d���"9s��?)Z�~B�Uvϟ�N�6��	�&��2�w���v�r�/��*�9�X#�&r=Th.l��8D�,]�d���y6X�֢�Gu��T�ȁ�H� ��ʯ�p�"���)�Y�^�j�^�.j���st��o�	De���S�������4�mVr�.�B4������N.�=�Uu�ߛ�����k�`�6��? ��uD�P�j���B�em��.�T�3b�ghIRjv��n00�
��wH#��i��s �Q�j?k��%�V�(�����#Qtm��ǝE�W-�4��JETĎ�ϼ���Vg�Y1ί_G@����Yml#^9e�3oT�c�
2�Ł,�����J;9�3�hE�] 9wO�~���f�*s�b������<�W�����ͦ���~��

�d5V�E�iv�hme%�	fP�"pe�|��gqŶu�E���>��Q]E�$����Gn��BaV��� ��R�6���ry"b�%�yl �P�t�-/sD�:;۽"7�ZX����Yj�k1�����4*�T"M��P�wZ� K�b�\�j]��!aΈ�ð�Ŕ�*��a?������~<<_rdPN���K+d��"X���Om��-��?9���ӹǛ%(We��9;Q/����DR^�Ŗo�*�i}5�U����|��H��o~�P>��5r��j���X�`�gzX�X����{?�����#���w�J���h������z�c��}�n�{\s�B�t&�Cs:����j�3�'i���)dA�o|�0����GDaM�'�>R���l�M��̉�[^�j��8#M:9�T�����P�Dٝ�>����#����{�!0?�bv:z���(��3p���X�kR��E��ww0w���G0ݠ���z?c�|냜q1�h 4�66T���#Ng�A��l	�u�ϒ���>��`䂆/'�%����t�k�����3�=�ޅd�=��4׸>���6kP��
��}�y�n�g�g���0w�0�{�}�I
�����XX[J��J|i�c�=�SI�O�ђD����^��k$`o%i���'�<�(*-_W��K��� y��aE�������9�?'[��NF�$�A�J��*eB� K��x%�>�y���msP|:yǁ��૥��f)1��>�~�c�i�^�ت&���	ϫg�Az)�v-�@��T�Ydz���<C� IFW�[��䠵R�%���\����i��߭I�/7a��PH|����]���g;J��T6�t�O�n'��"��/E����>�Xճ%'r�i|7�|��_Y4���PT�%nc��
���S>,�C챩bM�L������@Õ}�eM�/�i>��%�$ �3}�#��o�m$5�����<9��9ڱΞ���S��M��^��]����*,%i��vs ���~g,  9�����f�b�b	{�٫�"�E,b����[�R� :U�ٺ�疯o�9�H�����N�S!�T�w�����W���>&����w|��Sd��Ծ8��Mc��l-
��
� �%2�WY�ygb�T#*�0��l�{8�G`��H̑���3$����
`��2�<���z*�+� 䂓 P��ް/?��btJ2�	������.�"�ڀ�bҬ(��4�m��F��d3�Cy?�j�NF�f��O��Q-ЛZ�}B�#��L���޼
�5�i#n}�҆�:�CښPh���ȣ�L�|\��:��(�Jv�[Z���g��v��)c:xiy�,>��<6�W�P�$Gp�B�(Uu���/�ǧ�XOe׸�af�O��6������k.
��}
Ծa�\=�pL*�����=1W:������$D�ʣ/lxr��nk�����'�yhs/O
]�[��ޭȤ�E�Pw��i�}�/�1��_�0��0�U>{��@V�8�l:�s��M��?<���H��B'w��&3��HĢ�w:�m2�t��u����L�Ibn��3[�gKy�����:9H�%@� �Mo�/9�s�L-Q��ܙ�T�J�=J���8�}�}��T�����'_H�Iu�RB�����}>4� ���D+pG'�2�	��yR� hQ�������x�g�I��#؈j�` o�����y�4�,w��������Uin��� �1{����"��/��%�@f��|�_�N�҃�;��g��|�G>�8>���C,�����7����\�S�	��Qi^v�[�ۯ|��lu��,��n'N��T����f��f���_�SaIĢG��ʖܑ�I��#�������SG��^�]r?��|��}�{�
]�����s�z��%(��/Z�ο�mݴl�JӮ��y,BZM�|�����k�����O~Y�}�ĥ|���E���ј"->�Ҧ�m��)l���,���?7#b����]��'�h}�~���{AqmNB�x�_bҤ*O��?�Lp����NV�}_�{�(����r��dȜ��џU$�gvg�nڏq�Ѿ�퓲���xji��u���	qYA ��3���X�����;��^Q��>� 	:h��Y�Q���Q3��b���Ё��NI�rIx;�EX��g���+�0v��~���}���,�5CL�;���?[ �Ҧ�m9�>��8�A핞�7N�oR����z� FXK\f4[���l��u5��3�T2n�c1�!������įDwE��Y6�"!h��-<q����#9��{�j��Z���$t����!��օճv_*}Y����'M��X�L��WS�����
kB�A1�7H����9:6�bW�<�o"h��CN6_�y�=ZH�k"��vG��R��v8�]W\;z�Z�U��ǩ��7��&Χ�'J�$��\�\z2Z����6�+���L��G���6��f��C�DY��R�?{��,r
�`K��a,�V��b"�S	?��+�-�+k�� [3ȸ���������,[���u�7rЗ�8|V�����{���r�o����W��Y͜���X2�����%�uG&i)ԙ���B���R	>�|��4e�T]�B4w�q 9��lX
KL��G���
_���e�r�8'tU�Hye�o�ZDWz��h��v ֑x����	��>�i�X�@#��&�J�+K���r���a�<#����J Z��Z��JX�k�*�}�&������dnr`��;K�52���ƺ):���˛|��.LuJ��u�Uz#�M��=�cڹR���L�Tx-�O�~���|#; KA�"?��
��^L���3��L�f`�]dy�L{�M
6��v$��H`��BE�f������H.T��L��ݚ��c�奨Xp����.1ќ-�l#�	DX[�_�w%�K��"��|s20�~I�(m��v���������h�����^!#2�*Y�V� #�3���H������c<~���	��Ġep�)/DKRr����Y
k �=+J�J�t���[�h.wH{������	ͮ�e!����-�U�L��Ż�ݞ kP�eޚ��fYe��.�"���O��XFv�����L7�A�lC\����H�����-��O��+Me�� ����rN�g�¤��N�;��$o�˚`�R�Tʎ\��:�����iO�}�w��+Ow\�T^�D8r��֬�9�_�u��Ӵ��p� ����ך�]�Ybs�H��s��U����~���lg,q�ʣeZ�%}��W�1a[+Z�A���Z����)���f��iQ�R˻��v��'*���r,ؤo�5�Z������k;"M��X��e�U0K1�>��|HNĬ�3�^G�3��[�5��1��ŉOP��e�}���7��5~X�lI�3�Y����X��$ʡ��]s��la��`���W�d�0���&"w�Mv�wI��p;a��+��1�����97�s�iu'!�Y ����.ñS��������fQ��	+H(�O:�?�Ӱ���B{���]. 9?�y�!L�l��jK�pɗ%�P@���������6���KU6�s�?���,��9+]qi�]v7��Z6H�|��ǔZEz�S��jI������t�cRrԚ���|Ź�X��܀�h������*d+��Z��ʾ�(F`T���69�j��t\�A�!�E��T�[���'-T��\D�t���-/�&@9�̴`�^��V+���R�� �����Q���ƖP�?��b0��əb��;E����#
��Q9�G�e���O�K!-W�)�6L��%����������|+w�N����Jg�A�R	k}�}�hۃ!1
��b�,����O�sdE-O	Z9��h`�����Y��3b N:t�{����"&��j�78�[9~�_�o]� iG}��#�(�k�Y.^�%6��)��o�����fM��_����'����6����
�7�� ی)���"��K@�CSS3+�`ϕ;y�����k8��~կ�-��ꝊŅX��u&�˃�e�6�~�*`|�B�΋'���,�g���z"�v�X�$�O,�m���
s���pڏM�W7��ar�Aؠ������U�"����p5�bz�.�����"��r%XݮEK��-s��Ӯ�g���C?&�D��V�|!c����b�UP����I���f|h�孵1�����y񋸫�;��fM8��O�5�7Q&<�O��$%�;�z=Q�ez�p
���Q:.� ��:U;+	�Km=)D��9^�Q$����۹�Kr�8�	k�S��t��5�md�&�z��A��;�5�(TҳP$	�`#�6�J�n$�y�R�4|
�j���e$�8p����TQ�淌�?��D4��fw�޽TKV��|&�O�&9n߂eXO����$Uw��Pi_�T(�Ҿx�葖N8�[�}r�,����q����x�y��hA6���dЍ�_ћ�%WXe�'�����5��c��P��f�A�#RAR�L
�&
��#�(8x��Kم�J� 
��tk���(Op/W�11�j�g1���9�y�����Ac`�G���k8Z������ɂ�g
/��F�Y�������X0B6E�*ƣ��l�#�A��N�oY;W�cNn<Q��_m<%s�f7*z�T�3*��b8�SQ�o�A����.+SZJ���$�{�]i"�ͺ� �Xw�C�gF4Y��L�R�B�?��Pз��ի�Q�����"9x�.���;�����Eę�R�;���xM�v���@^�Z%Eg���\@"�scij����A�����]n�\�R˃�HE�,֙�;��Wޞ�sA�t�<�{��t�vh�[`]cu�����0$��w2p���_r"���~�3��@�A�8(��T N��-�7�v�>o��=�ZD�9@����H��?�r�J�p��c��b��Ə����������m�V�@�%:saz/�?��v��,�e����=O��ҾY�E�8�2������:��ވ�1����e;�<�&�]��k�g�j6k��o�Ȼ=Z��[�����ԫ(A1&�6Yv��_~���q��(q	����zl�/m�.b�'C��Ǯs�h��R���h.����+2��ߏ�<N�姈u6;����(Yc����)�dY������X�$��??��� �c%����Y$K�·Q�����0�y�}�y֞����l����+.8�G��حd3̎�aa{Xق�Qk����H��v���&��!�lK�h�7?ή������������ſC�G�܁�2I��H��h�pC 7��+��u�a�6xX��x2�m'Z���WC�O�H�V6�����z��@�)���������<�i ��9t�"c�zO|��-oVE΃v&^�|{�c������f7؜
����?8�տ|�o�
ؽ+c+61��l���{Q��$�l��Z�g�,B Y+=�X�N�a�>�x�TZ#w�2*�@����b�S�o'"V�{>S�������Q�ءZ!�9@w����x�*'�}�aMV}Y���8]6!���ŗ/��X����`�������]%��K�1�T�E 2r+���]Β�a�Є�x�]?�8*Dȥ�cw��
�J���X*�k�� �OE�wr`[�a���FE�Wx�g���5��FX(&Mw�r�&���t�
�?B�4��o8/���e�@�d�|��'���Rf� ����
JT��X�L.#6[���=���=�_�ìv�R���}IX�� 
)G`:0��/+a����\鷈�R���y��D�@Q�81�n�_N�cp�g{,d�Zᩐ�>Q�+	���C�;f��~�-#ώ?xN���} _�˱R�~`��:�7��bFg�v�B��
f��'Cᑦk1�k>�!�v|x�l(�T'���Q�L����N�����*��d�xq��ɿ+����U�1F�\��m~�P�=�ڗ�?��w+ "�ޓ�����R��"�j*K�[@���#�^afgXΛ�Lb��h^ܰf��� r����R�&"_��a����)��JGk�&��d��g��u�I����@�r|nRa�@e Wu",�k�������$O^�ڮ���Û�u�Y&&Y��I@���b;���c�R�h��y��>�~�P��2��v[�Td����ѷ2#�M�*
���P�����UϗY�kʛ�k��8��u�{m�~$g�r��T`g�ѭI.�@��_��'�Iz̼#$�@:�5J���/)i�Q�e�.�司{�s��<:��XN�� -�߬����$o���M����mN����~S���'�&H�{$����pG���x.a�DI�F SbN��{uy�C#�Ng��dJ����3ɂ^�.JݰEv,,�b�<}NTjֿ[a_`�%,���&�3�:�����*�Y���@�_�i�ݺ�&sN#�1"����kq����H�&�mA��Z;�vU?���}�>(K�ڻ,M6i�����iKߐw��e�,`��i�|���1�F051} 7�g z�?O{E�����M��]������r���͘ҹ�~�9�H(l��2q��8��|��������@�t�g"S�dm���Gз�r�w�z�X��*�q�v�/�#��%Ȼ���L�Q�v�>֧������ t��c,.�gA�}Ȏx�ލ�uJ�{�W��U��a��/��W���$td:?��#��:e��1f�r��ؑ#�u[�GK����v�*�d�Ĕ)I�B�>W|p�/2:.W�{�u��2��8�H���v���:��-H��B��������I����x�(!�
:LA��z�>��<�e���&�s��������� �l�a�'nM�ܬj�W�5�	�	@B�Bz~��;��C#�8�J��YD[�*�W$���������0\�ή�m�#
Qd'���P��t�[K��_)�N�%�1��O�PZ��� HsEQ�#��'|ҳ�t�����u�@����t�[[�F�M��;�(�:y����Ԃh�S��KS��������Lj��[s�+/ ��"����5"� �n��\4�?_���hԑ��2�+�WMW��wW��;�yk�aRz�y�%W�t}�F�n4?�PT'�a��k�*�E����j�'�O�I�!1��@�xeQ~�Y���&FR�P�ϓ�cC���]�')������������!�5���c�5\���y(�k{��;$�NCl��u����#�Жp��dA��0>m���#�ۿ�D(����R�	l�bIZ�Y�?��h��l�מ��N�F�S�w�!P��sgλ���I�������
z��P����������B���[��$�*��RfOo�$vO4s�d�{��[�L���}R>�X�����{!��k�{�#��4�Y���Y���/���eVs�"��⣧�P�u�bs[��͇��j��Gn���#��DC��y���!�y�aH����hJ�L�r�h�1u��,r8K�UD���!�)�w��X����l��B>��1�u+A��D����N�$���Φ�3���bSt�x�p)�z:G�;7_�䋫�i�}�J��=�WV��ڣa��5!�Q�7R�Y���JX���S���Vux��-B�n�L)�.?'lՐ����XQo��ЩRߙ��p�/`���3܂)lPp��	4����q�S��L�
�/�T���O�.��P��Gʂ���
(�]�ϹO_*f����F)���Johԯ����xb��n!w`A�N�R�XlX��F|��5u��:X@��E*���0E�U�$�T[��>o�ԝC�	���_�� fN��r:=�ƎrWГ�(*:�V�~�ϱ�Z�T5�T�
��~q&I���ؿ�a�M�ޚ	 �(�������?�+k�B��<���jG9z���]�'4�:�e�$�ⶱ+FwT������$�-d*#��D�X�R)!��C��rC��I/h ��;*�f�ۨἙ@��Zfr-˶zFH�H������S�P�4�}�xc��[@��:fg�zU�-�爏��P�&}崼3N]���y&ҭӷ�i�?F],_0��Q]�o�؍�/5x!b�u���S�ς���׎fOE$.�?��~�]�ӑ�߯[/�S>-I |l�����_j���pͲ� ��4���#�T��3.�9�9_��@�/�i��{x2:�5���p���c z���Ѕ�l{^7,4���z�v��J�in*y�A�ǈl��d����֕�}i���㍆ϐU�
*{��z��`iK9
�m�o�Z�ą�fs�W����E��������x����S
�yһSV[)S:�M� =$����<���L���Z�r���dg��b(�U����ڞ��٭ܝ_yo+��b|(�ܛ�QUfu�������JN�`�gqFm���Jzv�7��n}���K-4X�Z��6c>0+64���Ҍ~Y!��s�tb�	�L���#�y7�(wD�y�8���sYLy��+�J+r�.2io�
��-\n�h�i����T����M���*��+Q�Að�WP�V��&�si؋6�3�AbrTRbFlGE˫�-�s*<�z�)g;L��Mv\؛�ARP"�	�{�,?��v�>�ɶ
g����y�;$G9�r�����D�'\��ә�Uz��L!����r?Z��;,Cs�.�q�Q���ۊs���
?~���A�}]�F�y\)����L�٭�����B@?�^����w�t$L�Iu#�����������0�������
Je���8�8��$�N`���D��Ū�å��K.�w/�T{��K/�S��&^�\_��圿:M�8��ԩ
.�j5c<���7��,���ދs�ro��7��3<���]�' ������dCb�&}�R�۩`�?�HKP��x�A*"��HS��Ty_��o��8xw1/�p9��M&}\Lj����{
�m�Q�l��,��A�C�\��ᗈ/�Q��	��<������T���e�Y���6N�d`<��u˼�i�~�����b�l��2l8�����PTb���քxk0���LSsarS���Y|Bk�W�a>��F�|w��� 1���qS������߭ZG��G�F-U0�V��Ń�l���ùX��K�Ҵ��Eq%V:���jߧ����+>�@���{���IϤ;N�_��G?��x��ԟm�NJf��I<�� 5˯�e�~���������>�;�?��I�q�����H�"J_�Ł��vގ��ſ~�r���X"����w�0������ºe^�A9Uݲ�a�w9�Q�K�br~jD�~�Q����v\��d�˪���t�F}��+�c��\�|)�Ŷ���f����|�����Q8�TO"���I|�p�<��G����H�E
:&���&��?�^U8�O�z^�9>�>M��Nv�u�e�=K��(SH���5d�p:6_�v i�O^���X,A�baIj�b�g�?���ө�<'t��L�H/K��(��' :E����7v%�+��ܘunPYr�~6kq�ᢿIݷb��{vj�>�6���Xllw�A��� �m쎠��GM_'��?�_?���{]g_������+	�u���0����	$�zSiA�	��X�`�sYX+�ǯs�Ϥ~ w��a^��<�I�%�p��7��Yi#MS��$k��ޗ��5���?�����n;a2�111qc���#9s(���;;��%f]jW ���ܥ����e�|����>�f��]�S�Į���N8>*�����y��4��>2�I3�Q~O)P+.�P����%
�E?����ӵ�"� ߗ�,��g~N�uq,D�?'�m�Tnl3Y5G'��o].�j����w�b.G�fҖ�����çm@���P������ӡ��{N@��[eMM�Bڎ^�,��3����]���·e*|�s^#e^�m(e����"���"]T_wz�4[�L�܁���߈+D�<#���x�H9�4��:���$|����ݳ�Ҹ�<��o3O��K�E�ۍ1[f��g��Z�&oTnϸ<�T��cU���N�W�x���J���8V
'בQb<nV7c��lfKLm��{Ă��F��V���'�͞��W�O�oI�Rԓn�$��5���ӞFY�>��	��y2��d5c����b=��s�]E��e���������byY屮a�4���6P��%ft =�){b *�_��:{�⭣]����U�C^�͇��$=r�Ҋ�8ïKvCr���{�c�>oɔX���n�U]�ý;+�m@J�5k,D�N>uylJM�O�칹a��,omÑm�����Ny��J��K����y���`�`�.�埽\D�+t1��A�Et���rp%?��l��Eb��/�n���tT2�-���`5�^A��S)'��V�"�)�;�h,�İ/��6N �7.�,!��,n���GF�)�&��>��W��t����';�A~�}��o�Q�ƽ��3����D0�W.�ADBr� Q��r��aQßƳA�J_���`D�Bۙ��ჲ ?ηo��%�3'�?	%%G9��q���=�Hăf�#Tߺ068b�[I��n�#��	�\�D'.�9X$��cݸG�p�����(:vsʞ���y!�*m,:���z�=�A�V�f�FR(i�q��o�t�6������,����PU�֗�ϐ@A<~~�S=&`9?��_���^Qn"p���h-RD͑A�����Y��c�4�kק���oA��;��E��f|q�0�i�!���6����?�h�I�Kе����[���6��X�6���%g�r�Pv��j�^B���C����@�R��B[+N����3�n��J� �:�%��ӭ���oor������B�c�Rs���0N�V*� k��^�za��v����D�t�>��	�9N�,`���K� �&�$���5G��hH�#���'K��2�����@��3+P�p���y�e����(v,��o�_���¾���r+��/��X1W�#j��j�>��k�-Q��)��1�N�y�aA_���:�m�>���׭(b�B�E�ܰs�9����W���n�=���n�V�lg��!��yeq0�����hrZs���_b��ba-�guJ�wF�Pq��W�r`Ǫ�FB�(��������<��g���� ���dU$����c������u��;��u��JR��M�w�fCA�]�2�B:hӼ��V���g�N��2C!�S6��R��rz�݇�6/��L��s^�
T:�t��q�TC�/����4�8�ɷ�#	�{ycY�L�ܴʵ���B�o%=�x����y�a�_�gVz�	{��Jq�&��76%Au��Γe�f��*y��+J����ޛ�C�v��/�R��"k�v$!�v�J��mT��'�蝢��(E��}�d�:�Pc�f�f,�;�K����������������s�s��s�s��^���_���J�����I��ƴ�:z�U����7�����q���!m0D��ݮ�蒖��c�m+����-��7+��1�+u[/R"���7?J��9����������r�L7YU���iV3��(9
{���eK4	ӑ;�j[�@���gÖ��}����Ӛ�E�]j����Ұ���<�-<��w�p'�$���	���cac#c���x)ϣv5+�O]jf�X4N;0�8���29�۲���ڰᤥ�y�,%�S7<��M�xX6��s�1ګ|������I��שּ������W�����ː�&��r�]#^FIjGc���s
����uι��׿�Ե���Xf�����s�d4wE��g����U���1�����~�~�yc�9�W���skKNn���2c�pu%�c1�N�HA��s?o��c��3�*�m�z�ޕd�3�,��#�n���>��[��[��b8?z��3�ĉ\w������_l�.f<O�g���B�/|���M��۩���췍������ٺD�ܗ!	�{j� �ӫ6�Q�NML�9�_�Wr�*�f�is�I�����]��D�U[qf2h7��c�"���@��J:>yCx�`����9�/����.�w��pS`�>�G����`b�C'6�W���;�^�E�Z-VY̭�w��JF	=���9��\�`�]���'��5έZ�~A�����_�T�|��o���˿�[9��f��+�T.�M�y�^���%�mj:�����cOC=*�<4hǚ3���b�K������������ ��g�W?�ѬΝZZ��(�)����"�o�-K�W_G���b�鷞�O-�>%��n_O.��y��.�ѝ5}=+u�y^�/s;�d���˸ysv�Ȝ�7G�G�W���S/�d
b�����oR|��Zj�m��9���+��:|�Q:-7����_H�-lq��~]�ċ�W�_y$e�L�ڜ�Q\�Fx�=J}z�zۅ��� c��Su'
5����7_�q/������>/�� �
�L~�O��V|/��I�umEՎq�1Z���|;kM/Znuk_ؘ��R���Tt��|���<a/LF=g�����0ۻw^�1��>���mҾMR;�ʙ���q�C��Y�22�a�̤ꋓ2����Եl�]U�X���=Mʜ�EnSq-%�Ѷ���%�_�yP��~p�h-�zF���
�Lb��N��	|�n��^�l×xb_�I��;���خGR��_;��m�2կ�%,f�i���{����ޭ��n�������օ6��cY��2L&J��!�}���i<8T�M�΋<ZDiu�$�Jo�k�)`�._����ܥ;l�n�OK[��)�O7��X�g�����D�c%
��Ԕ�{
Wg���UZ�՞�zc���W#{�9�ch�������?��s��L�֙z����C�����<�ff��u~������|�$Ffc �hڴ/�u����P�z�&֟�m(���)��9ɛ�ǧ�Ǉ�J7*S�+ޅ݋�h�­��g���Ͻ�e{�BOY:^�%�D�4Pƽ��N��}�1_��r޴�X����E���*�u�D���&_,�w%s2F�G�:�:�ޏ�V�H�+髟�[5��>|e���dw�Aj��)�8�[�|�O����~�����,+~�7Q$���/0�
Ͷvb0Z�F��cV�ݯ������ӭ�~��Ԉ?�on��B}��i�d\�r�s�q�}�E%�i����4��Gj����W]���[Bw�����b����D8�a!��5�v��w�V�#��hˀ���}:.Ǘ���Ɔ^U���4�J�}˽�.��)�y\�@�\����p�(F�1ổό�ֿ�e>V>0����4��묤�y��d������O�υ�=
�>q���zR�5��nP��zV��۝h7���S	�}�KD�)�ǧN��#.\4DT������;�m���|[�@�O��f�ǋ
�{S������?�A��xr�u�I���~��Ĩ8�����p�۾�z��и�b�X��l-|�}T�Jyf�\�(��[�"v�R�vD>�~I�H���x�k�<�$�PT�kB{\M���B�]�N{�9]5oiRR���YY?�a>^#���QL^�N�'M[�E]���:�:�g�����6^oZ�r�y�'b��aY��s�.�X4�,}���ihbK��w��y+��n|�>ʵe#�ofO���&�a��ΰ{��>h �L�>�>	E�w���n�9���6{�
�o�3�x�L.��wv����7GDb�]�z�a��n�h��3-���΄x���.�/�ʳ��jVa[X�.�<�,&�q�	����M�s�{���s�aq��a���}Q�O*6	��n`���T�d��5 ���WeW�
�	�<��{�����ۻ���g��Q�y��p�������[��[��7�3�G�_��Q�*��;�P��_���z�s��g�C��E)Z�Q�o8�J��eS~�Z1��o�Ck��n�NML�ۅ��v��]�d�_y;��6�SnI�A��7J��K�Cj��1��sԖ�|.��Yb�y5�"߃��__�ל������O��Ӊ�R�#�E��Ϋ�ʧ�������i�ī��e܎7�b��Mc�h�����myg�6�7��hR�D�,l�^�����S�l"��j�_�ϳ+����&xwj�g�v����ô?am(�`��	�]�񦀐�}������ߺ݇
]�M�����ɠ�h���g��O�8��+�?s�z�ݪ��9�ߪE\��w)��9c�7�0��ϟP	�O_�i��ƣK$o'^xh�S���P�zN֮�|o��.̒ߥxw��y�\�%d�i�H��/و��G����g�6?6�b�.SYO'����wj����+r���=�<�홱�K�-�Q�O���s8Ɍ����Q�cKʳ`�Nx$�g����������U��#c6�������ʡ[����v�K{L��)��Mt=���܆����$���ك0Ҫ�����j�ɟ\�;+s�b�SG/
�,��mU���V`Wf�������>_�x���iv�.���_{�V��Hm�K>����j�qS�����+冋�4t��t+�Ժed:�w��hy!g�'l��JÎ��.v|���wb�/N��11�q֊����=�Q�6��o�vM������ҷ{������&q��^q�iDA�8a^��>�������և�*W���I�T��k袘��Ч�,l������Rڷ9����i�&����wO�ND}r�{>g�9z�i���b��D|Xe��J�7�=:��/jlx��!y�x���r���=�7�YR����/(�������������\��ϧ'�vPW�����=ee�t�x����i�~�-&��&��(��/�p������ZZ���9���a؋�k�Ԣ��͙뿽��4/��h,��\������'���VR�Q{/��Z�IJ��Ms��;.��^�)ǋ�>���c����g��]5�ʯ��L�c�U�>�j��iv<P)��_;QW�n�?�պ��n���%G�I׾���r�iK i�����}/VR���C%�:s/����x��1g	������ôiK�h�/�����oJ����)�X�9:u�{u-v��pF�s�{Ea�7Ocٚ�9>��M������]y�8a0��#L�hʱ�o����NOQ'o��.�����S�z&P�~�2]���l}��F>��,��:��S�W�7�U���u�V�@{!l������_6C�+z��<�V�UⰧVR���h��ܫJ�B��ˏ4�q���|0�m�aȾ�ݦY�Ǆ��)��~sNȸk�(s�Yu���+���z,�]���|8m5K{�H��Z+j<C��9���n���{<M�X��>���Ǭ�W?)in��]���&�w�'G�e��äx���;�rb���!;�,�{=l����}�@�\�IW7�}��㇬�����F�����SҿL?�n�5uַG���uu]mZb��.M�9��T�zj�f'9�^4����B���P�/��x�����I���n�@ �Ǒ N�2�3iM�]}��l�UM�*q�Bڇ��ENF�:�{��o[�-m�j�j�~D��l�fzJ ��鋧~�+Z"���wv����w��j�7�#� :�~�a�Ah��i����D�+n^��Cw�Y֩�����u���xmh��[�D�o_�ft��H����J��P�X�D���!�~;����Ry��{����M���ڔ����'��G<�Y%�?nlZsm�Z�'�\�j���{�Тڏg��Ҏ���W�?nM��ˇ���yn��6U�vEF�B����^���T��?*�>ǣ�&Ls��D��ģ��'��`j2���g�j-N��u�z�\^l��+�0Jk�����n���k&���7����T>/����k�e�m,k��*�a\�^�w�~��yo�%�Fn�K��{��e�<N�%��O�V4��n?�\e�d����P�=��6i�>��,ǔ���#���~>��{�ޕS�#�G�G�)sJiM�m�վ�����ΩՁ�Z7�Y]i|?��v���}oXaY�9y��O���u�7�m%"9�G�����<��ϧ�N+��t�MN,ʌ������_��#n<��l��N1�l�ٱ=p��*OK.�8I�y�$U#��N�<�ױf�i��*��oy\�5M�s	�~<]�){\�t�S�C5�uO�U����㭀���C�yJ���������A�+�ۄ��=,�_�r8e�v����q��Z��o�y��V���r$wqװ�j�q�'��,�\T�I��\X�l�|Fv���ւ�L��.���z�Zb�r�Q
ơ�g�m��nX���9�r����m�����+�]
U�t��xS!�v���y�g5/*��ٟI��yɹ�|܇zi,+�'V��q�}�e�Pv��f,����,��`�Sj�m����;>7�~c���MYⷹM��~�(��z�������s����S��j{P`e�ʛ��)G���0��=\I����"~3�n<b݌�3�L�tL�*	��T��������z��\]W�<�(�����^�������?�:���xH�P�u�T�V�*�oK6��T`#u���̭�:�m���h�]9�X�aE:/q��F�grL-��4яK����'X~�����䕯�+$j�~�<PV`S�z�巀߀�E��N�\�a�g{&I�_�ϻWǗxui�L��g��Jq0S����l�!*+<9D�UK#�B:pz�����}�v�ҿ�<�:�3�c����"��e��p������_Yx���XK߮�����g��iK�?����Z1<��[uQz����Α�ŏ�kK��iO/W���ݷhI��v��gf+7�T�d@��	�~��4oQp�e����E�n��Gm�U�X��Y������d=m���✞�V"�QV���νg]@X���Uz��Zr�)[��)�ȁ�h�f�C��.-�m߼8Y�k΃K_%�ww�"�'�~�p�d��C"�b��зCw����*��/b���w�Y6�����V�S�g�X�0�حԾ�*w�����W��H<U�#��wa�;C�`����s9�F_C��za�����n�O�}�p�V.�Ӕ(�T�YwC�?1�E��oV���9��+Q��48LZ0q�	��֓�U���#�G]w����*�׾G&X"���󔉏Q�0h�Y��S8�A:����TT�ٷ��<x���C�o�o=�}��C5�SQ��9P��=	��*_�<;r���˸�����j�+àw>��+�vh�?V��Sn�>���<�\0��9����u��EI��}=^�=�cѣ��︝y�?٢|��`���w%lҤ��N�����,�A
۵$n�݌��94�-qx�S5�p�BՂ�\��&���W�`�Ȗ�m\���zk�M��O����}�D���o���Q\wZ#�];'��8��p������V0�z��{U�Ò���
F<Vڻ��m�݋_*'2߯#�1WB	�%_䵙��׾DX��>vŻ%w����q.�J�Ej<6@��y㺮*˛~���^�#�x��-凛�{�3Ft�ɒ]�^.�崙V�e�IR:Ń�Ld�:<�j�ߦ��r�U7�!�պ�J�asS�q��7��?�xb���Dq������o?����݂�'ory��܊�6r�I�%k4ɍ�D�x�MA~��������_a��d���ݝ9��5�򫬞��c�����t��^�Ԏy۵�ڪ�:���H�Մzm����5]r�C�X����|]X����;<��>+������ɟ�*����Z��Y@kJP?2x����Y��2�����,J:�� �:��?�t`*-��Ӕl]�azG�`[��K�&M���t��X����O��͡��ބ��=J��_rM���FUKb�N-���?�T�`?YW���)p1Xb�?c�ܟ3,���g������W�NW�j�M��'�.^f*(�w^�?���XU���k~�)�o-�ǎ��1,O��1�ʛ"�b���c2�Q:[r�{�h��_�"+�}Mјؘq&Mc��-�a�kQ��N�[���bsE*��o'������|֦�=Uje��S��8�����his����֕�W*J�
�jj�z�~��d�%t�6���EG7`�<���&�.��bYLx2g�{ұ]�:��/������7)P~25�Y��u�����I�������;�gH�z4���"~�s���?�jv>��#��G���n4m�xt��������\�+ϥ�9O�~�kH��>��ٴ���O�5��怟Ϲ�Jκ�C��E�(o��mO�p�b����V�<q����?�����F�%��.�U{6�-j��{�r�M��VEo��{���-k�)ɿ<����[>s��T����x}x��B�BE��&����oW����\-���l�C�j�{�0�],{Q�&���%\�Z	�d�Hϕ6�n'�難�MJ��!R�/ރj\ZgI���.�s����s�m#+�O��7~�i9��c���h�/�d�E�CԆ�^D���N��i�ɋ��8�~��7����\W���7�\��b<�Xy��
N�v����מ3�A�u>�Z�ɣ
�����)0��,=h/ꜻ㜤�ܛ��~��-���:H�a���1�[L9��;����pFzK�c�=���J~S'��q��b\�M>Ƿi_i��&��^���R��� �*��yi��F��Ãu��i#6�Y�����l�=�frTQ��;�\�!x�/`��'�؉;?�o����F2��W�f���d}߅�;���&u�|J��RL��'�|���N�k�kT�H��5V�B��o���{b���k�+� ]Wqo._q�<�ڻ��Zb�O^72��S�-B�^h��3aRV�|u����ʊAOxP��S�4y��b�L�"�l����e��#�w�f�O��xq����hJ���I��}�o���]�� 	�D?���s�;�OZ<L�~�W����+�A�ІҪ���v\[���=��4�Kw�i\>Ns�o��yi�k.@ӺO��0�F��=�t�E���Bs��q��OMmi:Z/�ۥ��g��k��S�_L4�|�L^��k<�"��r0�͡����$�P����H�.��&����x����J��-YS�}�m�5.U�K�	Y2�D���K���/�W<�������o��
��{gB|�$I<�?Ё�S�3��[����Q�ɱ<����]�k!�1s�c׮)�u��x|&���&�u�V��s3�&6��L�5�q���#�f�ՉG;"�]�w�T���M�q٘�>�w�H��k���]wr����CVO�>~>����.��K{�2��X�����N�>��n{Ɔ����r�Ǹ{z�a�4:���*	���)��&��&��Ð������h���Ӌ����R����oL��?����1-WC��rW`�O�Fs-��7׾�<�H����r���8�|N6��vO[ p
(䍄�K�pD�*��;�n���\������3�vefO��n*�����蚉$�49v�t�d�c���Ѻ����[��������<xpN7�X�/V���[(C#T��ڏ�n���L��е��Ѱ�\!�R�B瘽v�l�&�����w�Z1���Jo����菻����%��_�'E��S��	����[��(�*�V��5g�IP���y��&/��W��)�n;���e�o����m�"5_$T_K�?�k��wd�½w�^��;v�����.<Z��Y����M�+��l&q��K?a{7�kR��:����Y��1�I�B��W�_�헒W����Lm;3�>f��n���wK}���KJl���Y���)[��OM���s�2����ύ9%p�����s1�s�0+WVVn��e#V��8�K�Ju�Q�}뽂�jw.[,��>�l�΋!�:&����ȏ��fq�CAwf5?�$��شcC�≟��޶`o'�:��6�����P��/���h,&�Z �5��K�h���xʌ�]�񂥼��o��<{*���JF�A���鈸3R��0���0F9��fDzi����T��1mo�,E�*�B����b�^Y�n��D����{�`�8��'��cq�R�)9!�ܴ��/���T,�����Qj����q�z��1J:���ȋ�M��Kz�J��MZF�b����J-5�?�M�3#E�1��<������SW���ˬ��W�Ͻ:\5�9�����k�W�t���f���kxTv}Kh
���1��������1�|sB�U��I	�ʋ[�4e��܍����ȍ������,��ӵ�J����X��0 �Pvq��阃���ƈ["zx���s��n�\�y�']u���P��I�q��;����L�(����ٙNK�C;צ�S���\*�x��ZX�����R����������$N�+���M9�k=���x�'�w3Ft
���Y�Z�ex���:�E��F3o7Dϵ�0�Aܥ�����I�z��_?��1ʞ����.�+��.⣅.�)�N�n+#.n�k�,�@㾯�όj��PFTdh��0������e���u�bo�3ք���u�1b�GtX�i��e!ACؠkP��H8k���� 
y}xb]����`���,��fj4���=u ~�#
�O���X^�P�d�F�.8_�{u�Y�������~��t��"�#SA��IvF����X�kӛ�����v�e���<�j�ؖ�(���1�4?�����Ώ}L�"�-��M�<�zW@67'n�}c»����)=��*iکup�x�:')�)�I��3Η�J�	���a���%*-#�5|u����K���
�,�.�Fë���;�0킮o5n�c������|d���=˓t�!��?��|4=��d5T�n�ƺ��V���5oL�FFds��fh,t�Do�_`�;Kk~�2zk��,�s���H���&o���u�Ē���Z��0'4|^�)H#%-܊wBesٳgy; � CA{���i�&�[�b��@�'��s���כ��|��=���ҏ�<e� V�ЧI���;���ٟ���t�3��$��J����l��n��j�0+��^ʈQ�>�2t+��$�J�#��CW��s_�� ��D!_����=J��Ҁܺ�+4�Fޙ��@�J0$ѫI_�)8�X[#���Ǩ��}1 }��d�p#�h�ff��s�}��I�*$��e�c�SO%7m�����l01N2A������涊m�sb�aa�D$����ey�?�4yH���N���?{�0�rDo��I0�m�vo�Լ�*���(���g��Q�#��W���܇�z�]�4��M��
�@|]��1�O�����ِ�جB�;0��L����HK�8k4�a6dh�� ��Ak�� |������ȳF�T�'�����Sv�����ќ�h*��]��Dl�m X��/	����k�1�ȁ�Fx���#�ťqi��q8C�hߧƤ\��^}*|q��D!#�?߇r�ء�ɇ�Ih5�۫��uS���т�U����az�BQ5T��S�6��o&!���?��x���>�9彣�Y]@>:��1iD*��Ԇ*;B� ^��E@o����s��t@+���=Ϫy�c�V�mձ
�a�ֆ���lH&nw�sr"GtΜ�����0�fD�q���X��vd@AJ�s���Bt��S�mD��[��*}O����e^����~d�� ��@|"bEY)��Wֻ����YnS*����|`1e���|r��z�6R���lj�W���8�Z��~���������X�s�<�{��:�p'����Ǆ|9�5�8�(�R��hG��?�^>�n�K@��{���G��� ~�T��+��)`�"Gr.�aj{�Ėd�i?}YiF4��:�}�ⶣ��!�[�f�}o�P(j�[oޜl��P(�P�3z�=�`ɢ	r2�]3��s�#Q1����\wv'JR��l{� f�Y	���b��/��O���wļ��j-�߳�l���٪3�@h�V��!�#橭V�>�Ě�}����=��6�Iy��ȉLZT�b�w�	A�ڣ��Î�x�IpP{,.�(����v&�=|8�-����X��J5=�퉡��6�n>�����5�ak��ຄFF��ng�=�����Mǭ�'��O%��)`��ec��|V��#�'I�b/�x��񷿞�'���D�"L��{{�'����lD�3����S�<vsߍ*�j��ԓu���(��ܩz��+U�C�?��P����폸u��G�޳]�JBv��H=8.����}�����S�A��9l>�D�<�w\-�t�#K���������"#��S\G��Z���=�u�d�r~lpI�����G�aO{��ͽ O���B	c���@��o�a�d�#��j��3f����}tƿ>vcVaVaVaVaVaVaVaVaVaVaVaVaVaVaVaV��z�?
����/V��V�.ۯ"1�A���^�;, ��w��k���:�ή���:�ή���:�ή���:�ή���:�ή�+Zw6D��(��t�|��~�vv�]g��uv�]g��uv�]�/\n���׻ �_�2�ή���:�ή���:�ή��6g^����\P�g�gbE�3驖I�Yh�&��-iJ�W�������*�MƼFtc�=v?�u��k����_���j}�bh����z�Mm|����l�g��+��mg��50k`����Y�f��50k`����Y��_P&ߘ��d���7���|K�<��-���(/'��v7���2:������wb�wI���|/����r�yc�
s0ڈ����	O�w:�������ʊɦ|^orDor���?���B���RxE|�]�,9�:1y���C�)F��0�ɸ��?��/��,��9o�FM��:i����i���~T��b�\#�{OﱱŒ%�e��'*����0�'>\ՈY)G=��-�H�X���I�*�������3T�W�| _��WQ�ĤFA��x�~�DRY����NL����jIc�b�Z؇�T���Pu�z�&����X��HN�b��е̠"dF�,*��r	>�� T�w���pib9��nvb��ɸ�_Ȱ2�����&����߅?oUC�,E�0����y��|�퉊
�󏼃%��Ɵ>��iQ�rE_��(h�ہ}����)�7���|P�F���`&Lp�rl6t�P;'I(���=�`�E%��~�O�����{)�X�](_�F��f���N�r��\��kޝ;1y'׼���2J�؜��ڠF�ܪ���&�a�np1�/ӡ�1"�
�n���'�Q��Ȱ�,M��l���Tx�(�����%��>���?�SL�u�eQ=g,�∽���qΑ��Q.��!���TB����.��$����'S��R@ċ�	�G�$� e�B��(���Xi��sl��w�nF HB��y3ԑY6�}9��t�O����g��%N�* Ჷ�s��n��#��+�3�#_~���>�3 F�#n�Cʼ��<�����]�[�!�`�𶙡0����%`�O�y�ϟ�d(#�5�9|r�)�3S�?��Kt�Iq���nHQ�*��ݽ	�������8TN37�D�!t�7����l���q��p��~Ri�yG9��Cԝ�I��2'�*(�Q������F�, "r��Vt^)�/���-�����QVe�ڂ���D��%ePbMr�T�2�&
/���$�d�Ex5�����L5z�ո�����Y���Ah���f(��iAI�1�t��oj�ā����/�d��#da�'Ya9C���`)�K'�Ā�5�#�QR�/��30
���L��ڸ��tP ��Ӝ�IBT(��)(���q��t\���ÖL�I����� D?�J5�K'�.�U>1�d��Qo\�+(�DdREPܷ�<Ce��U����� e�T�V� �ԮAҍ֙��.�+C�T���Du�#���w��2��əR�t�֔���݊	zc"lT�:�����b2Ȭ�����>��C��6�s��U �Np3�u�L���Qg')�ŏs����nO�Q ,�`41�H�5� "�5�Te�L���	FʕO'&?ч�>�\+} ���F�L-��"����F�́�-�ٱA�]��WPg�D�VC������98�﬎�B�Q����3G�w�,)Q;<4�ϟ��������IK�0lx�>s�l���������N��V&��57���!��&(7��L��upX�ߐ��d����q� ��>SC�zh��w�ߊ�0�3�^�A㜭35i��12��*]?�,7�����wa�S� q�Iy�3A�v^E�P�2m�;ᝉ3ѐ�
L��͠�z�D1p�DA_Tğ�NVf�Pј��)���qj?�r+���(Cqa?�\�.=�u�M8Ȕ����	���<�F?�PCE��qxp�L+�Mx���H�S*d$�q��������d�<.�a������o\
�#�`ɝ���qѡt����X3tdt�#�6@GF�؄7�#>�
N��J��������ѱ	�0i�DV��Б�R�<�����	�+�^�A;�� :��������ꭔ�V���̡k��Z�2����׆f�<8�C�����:�Q��@����q���KG�A�Aߔ=�L�+��S
�����F��[��鈎�@��}))�a������l�����«7�5���u�'�53t����Eo��a��T*}�����I�����|Vv;x�`�8������h�S�+g~P��4t�I-U��wH#g��ۣTj];Q��\D�}x9�H0��; mF[d���[r��	� �g� �� �_��'����n��4���.�1���H#_[Qa�1��G�Ժ���]zR!�E���O��U����Ol�~�K%B� �Q�����2�5h��-e	[�bOQ�����|�O��>�Z�'BI)·r8n�ՙe��4�_6T��Q���&�9�}����� ��^8&o�N3�������'P����g\���`hC%�}��%P�i3���@Q�l�5�m@ABܘ�����م�l�ɏT��Yd�@����cXLPv�#��CVW�2����d�eP��N�����f��pP�gtȍ�ƕ�����������"��YܸG?��ɹ��?C�S!��wg����J�C��-�h�5�!��yS*���U���ȡ�D����C>�T&���^- �&�V�7���'Ɠ����H	���ߐ�^�E>5¬5�v|�BD	Qb$n������/�|�Ռ��F�r�u'����\���F�y���7/����F�\�An�z����qo|*���$���+�9���������36;�ȫ���p�re_���:~R��D_������v�Ers*g�s����G�f��L�N�HS�D���wKQ�%�@���Ar`���ޕ��Gy�����r.�.B%��3ݐ��?�a?@�o�HmӝI%�t��oVָG��S��:@u���%�� �����$�c&MG����Q������g�~�x��b��"u����
 �9�34�T�r	�����3I߹&��1��b{��w�@��T�u�f��c��ȑ WVQ��19�}���)���:�|~/��;�zO,p�#����b$��޻�=`���zo�z������`��*��,���\4�^9�Q�G��Y�ȋ��1ȡ7�c�ģ�NTQ��,�s'�5h�(TU/�@(��J�	0灛{�I'~��M0|&+y�����>�N���O� ��0��Kj~W��$a�'�L�K;QY.���Uǰt�O �*��~ �W���Z��_3�F��@�x� Jsа8���%�Tu A�Y���p�ͽ�d�!���2Q6�}��d!��O�42@X"��M턽J ��d���s_S�׊��A(�(.�*�^&C6CR,�2l	#MG(]�@2_$�F�ޢA�Yr�0���.i� 4<��R�W�$�E�!+]ڎD_A�;�u��Y��h;��N2��:��]����J��!K����-c���"�!��%%�ˬ�;�ډ�o�{õG3$;2(�U�b?��$F�#�E*]r��fGجQ������߲�BBpݡ�f�:K�&� slD}3W�N�z+~�D~H����K��sI	��^���.)��ώNm�{��=��܈z����F!�A+�Cw*���fT^�p�3�	z%~|�	y���M�#ݸ�tIl+��c�� s����(�q����-�� �����qX'p�n�鉁��>�I؋d�H���2�e3���Jګ{=X-�[zs��Q���Y{AF�A�*�1��L؋���n{�,��{�\��ڤR/s=�HF2M$�YiSK6��#���{7�#{����"�˼{Af����D����Z���)G�"^����\�'��?��"������b��(�%��rȗA	!�B���U��2�f������-FSR3�w��@0#u&��9��߼�$6z��KfX
��RtĎu�&"�:��f�����tC��9�̇�v�._���X	-Qף;@�r'w�є�:Rż�Ԥ��"�	|9V(ƕ�(@��^��IG�a����8���蠨��h�$�1m!����=�����A,�B"D��Y,�l��� �1��/!�_���5��)���|��Y(ʖ����I�e������)�/q���;m���QO2�iY^�EV���r醌�`�����dt�T4���yg?�_��9�~��~k۝Qhs�P��Y�12Y�2w����b�e�a81;�)R�@syM�q0����G"� t�����5�B�`��cq�d3:j/�ƚj?B>4�e��C(��HbO�RC�E$��˭�' v��-*4,��"�hX�Pǰ�)u!��Fj�j;r��5h��f�Є�(C;Cmr���iY~oL0h�\I�����a=8}M�VDZ��Nk;�p�7�S���BC��Z������s�[�B�nPAִ��Kj�3=/���N��9��(�Ks �	���0I,�-u�Hڔ"��8@j������1@�����~b�0��Ajw�!���?>�f� ;��\N�I��H��U&��&�r���ć�*b�~�Xp���A8P����zp� ^,��	�p»Cd��^��l�����^���_��K��[�����(�}/�H#��؉~œ���!�~^*�sA��S��,h��\W"��,-��q�A}��Wd�w7��a3�ڋ׼$W��ari���� �]�"]��L���D��כX{H)��:N�"�.�T�;,sp
�&�#}j��R�Mkp���a/��Z�S�	8�pk�AMw
HW�2G�i8ő�5@J��"�ӹ�S@*����zrZ��7t�HqeM�c�^й(����C��q-CK�h��ʐ��A�l
~[��&4�cI��V�HQ2��6��؂�]d�w�.�V�܏��7�2ut�?��&n�e0���2�g|�B2%\c�[-#�B�3���yK���c���{�'��)�Ռ>؋dx�wܪ������\�^�7�} z�^3<��2�g~�B2�P�!e& W�h���$;���>f�}z�p=�!B�W`/��ؚa�2�fx�^Hw�M�w��e��^8Z*O�L�5��=��C�$��8��[K�z����G��K���83c_�l,A� �%���6���"��4���1hkt�}�YZ*�*��V�F,��%\Y�}�PH.idN&ƪj��&Q���Z>���A���~[ɕEe���s�K�, �����$�md�Ҙ�AÑ��Mn�NɅ�N�#�c��M��c������O����K"�2n�\ko2�[@�����������<#�!	�w��&A���B��&h�� ������jЂ�W��(m���DH!���@�f��3\�fn�� ��e˸�P'�=^� �N�8IL'�j{�n���B�A(�^�s��'!��pԗx���9u���{F��qV��X�c_���I�J��C,p����]�2��B%�b%Jˉ��:�-�F��������z���<Y繲Rz���	���1(R�~��bh�3zWAoٍ~0\���bYxy�37G@�&�b�߁�*
��r���pG�.�sWֳ�����y?��k�O�E��`?�w���rsą���%�2D�I�X
QO���|�C}���M5s*ʅ˭u0�|-�:�0R���ڶ:!�C}%I�R��\��-�6�ؑ^�+��g�Ok3K���:�D�#�B3��Ϲw�Y���y� �t���[��[qcB$��>f��������^�'ޮOQ_��<Q�80�E�o��Zd�+�<�́1�Hx®#�����a	0�+��a>ai-��E�p���a^�e��~^�m��0{ �2R���f��L�$���90!�Wq�4�V�K*��i�8�S���B�r��0�?�������p��'s:��ӾB�T%吡VѨ�-Λ�SH���:$��>�"�
�>������,�H"p�2��V�3��(R�/�G,����A2�~�xH�w����J�*��'���~��$����%��`j�^����
IR��]���� Yx�O`8d0�,��Ӛ���u��Fh8����\�k���[���Dϣ��W����-�㋨[�}�+Ε=_���D&Ae�!��	�P<!�'!<<�����܈��U{�m%����֒�� d8�_����|(��3�6E��[�Z;�3�Ǡ��!�>g8�{�nPc�!��N�A�((E)�f��j�sGw��!T�<<H�Kkĉ^uB��7�-u� ��Kg}QvE��f���X|�s�(�-<���_ο�w��";(�Γ:���҂���M��e~�/�
��{������J�Q���:g�l�5h-P��xi輦~��F��f���,��#^����rYZ^��يF�<nP�+;N�E�\��"���@��A��=UÀ�[e��F�z�3�B�mB 4�`@�g�A�N|C�*���ĩ8��,-s��-�K��{��b���rnD4%�4��@0��|�^��ږ(��
-nY�,�3q��XZ�H��e~ځ��f!W�g-#�>
�p=5�{E���-�ӎ�e�Ұ��~��g\O��'9� �����_-|/t�F���[8�p�p��,������O�$�U�����ވ��0x8�F�t���ކ��^gY���kv��/�!��B�����Ӗ�v�[H��Ar�vnD�h�!E���E�#B�=K+E��y����zrT����<�^g�ۜ��M� �G�F#���FYێ����Hb!}Ή]ڡ��tfs�3��K����D�Q��J�ڐ��(,�@JG_9�r��"r6j������@�1�"� ����#ކA�)�PGצٲ�e$���XQ��+��b�E��r[�sO��9��>�=�yϹ�f�n��R���:f���g�A8�3����Ƨw���s#$3B�N�_���Ƭҹ+�O�W���@<��� �2�* &�u���UR�w˅��Ư��B��)"�I?%��g��{͊��y�sʂy�CB׬�OȲv�ID��c�aD�����R�O\Ԥb���W�6�����S�^���g�z�=���E�B�7�j���a^�R���0p���M�WlQV��*�K�?o�>��{��^�g�
Y�Z?����9g��Ա ����-ɏLH1��A�WZ]n�M�8�=�]��0h��Xh\��
��3|D@n�o���u)�jd�i�������R�O�!��t����Ъc!j���'�-�x�ʜ?z�ڏ�46;��|<�������p��;tE��p���t���f�_����nu̖���+��u�ަ�cs����z���9���T�0�V����<g;b��V[Ƹ|Y��6�a��QY�$��x Qev-m4�h�,�@�q����S7!5��g-�7�h���̸���dÌ�cxo���`��|�]K�R����º��g�
l��3<�+�Sf2+bhU�Q�4�zݤ��+�_��u��Z���R�a\1H�����"RC��~	�R����ٰ\������^O�&$+n� �Ld�b\�,\ i��)5�J_����ŤtJM����f����P�{�\o�R2t#�e��ܪӆ��\y�a��];9��g�PK   �n'Y��T�Y  I�  /   images/d8e70382-63d2-4b8d-b385-7bc04a585f98.png�y4�{?�ʐJ�P:�Jd���̥m�����LQ�E�!6���YC��͔B3l���]�y���?����w=g���s��}}��s}��{���@GK��ɀ@ ��\���@����t�J��2��>�ˆıB�T1��LĞ	��(O��5Y+�shkK�s�N��?��O'O4��������?$!�&_�Wd��#�nm+�wQ�"
�O������������9�s.�v��edd�ED�EE�������'�W�كh�wUm<���]=�]�y����t��T���#�cm�gW/wGhk+aG'gO��������V�����6�a����\q�'� �v�S�����E{9z�+�D{ڸ��x9����ò�xX���	�V�'������no�g�sh���s ��hk2
"��������x�o���8���v�����j���g����ne�P��n�V:/./����K��W�%���V�R�BV�b6B���B�R�2Bh1	��b"hI�?��G�K��%�*!*!*)!s^������ȟg�����u/�[d����_��#Z���K����K�v�GB��e*9����ؿ�וLA/�[.���=<�����\��>P)�����]��@&���uGEU��7Z^�?/�����Ȁ
����T0E�0Ư��y	���D�_wYkً*�hMQmM��gd�ťEĤE �dĥeD�$�%�zʊ����IE��2E �^��r�7���6�Ǵ始��˻K�%7:Xh���yѪ�{1o�15�����ܦ~( ���Q�	j��C��LN^<}����ҩ�;�~:߆f+���#u��Y��N&���:��uS��|��=PiF�F�K�]>@���QA�@��A3×�O�B�������'�?�:j$��z�}e ��h�Bެ��5��좶�{%R�,_���Ja��ȴ�b��V�P�B�,�=��ʛ�,�[`z�}|�I&`[x�KN�ouL5���PѼ�������B��!az.^��@0����ܧ.���\ 1���gg��ݿw�f�/q��lĐ:�H�C�*�ds�s��v.����޶���v���'��p�����ǉ8�f���^�9�����ʿHX��u4���6���;_��)J����N�M�f*8�υZ�V��}�&xw���������;�+�z��(u��A�����Ԙ���<��i��DCI�����2���;�Jy�����9�q��5M��j�s#�w^T�o�j�&��T��͎����#�A!��ό��[�KQJ������3�Q�&�
*�֝%G�^��tRPB��x��j���K+T"��,�����2�X* �;�!H��T+\je�;Z�z���v�x�/m7$�����К95b*V�&�9\���:�v�u����ʴ��J�!f�NC�J��{1d+9c��I�r�L|��;k3�I��N5�@�&X�Z�����4���H��tu��*�V�`�c� 3䭀�P��z�W[��7��Mk��1U�C�~l�_:@���v�������q�`�?C+�{�{�Vkӝ�8��}�ТU��
�9[3�=�����(%���G ���z&8/ʣ�ڛf7R*�h�������F�ʜ��"�H��na���Bj����fmt���U���fL�`���z��N3��CH"k�͋{}^q��%����
^v{�u7���P�>BD�!!
Y4<�.O-�M�a~]Br��*�E�ކ<��L�7;,"�;��&l?��L����=���~�D�y�c�5e�܀@�Ԉ,xe�rfܙٍ����F����YKM	')+��R�����Gr&}W�w�B�
�׽,8Y���=�8����u�&�>����|/~��Y�O�@ ׊��s��G�.��x����r"Dh!�2WT������A@��[3�����_j�h,�`*<��&t�Bf\ TrB�NA������.�-קP��	�\��$�DG��Z����o/�-'g�3,��H��./&�nx �Y!��p��q�C�@�E����"iZ����E�	ڵ�t���~?H��1BI��Ã@H;S$�. �S�B�.]��n�������'�?����N�h���s�fU��N�9�o����տ����

R����,v��	
�
	���j�#��濋yqs���F�u����z
A��,�s��Z��������l�zsv��L�J:$����܆��,^�"BW�B�q���e��l��N�[\�������2�)StH�&�48�+���4}
�?Uf�)�.������l�+(�����=���V��-��ڕzs��nOu����H6M��F��㻒ع�����c�Q�MċT�qsIж�`�l�BbpFֆNM�u�t�\%b���lIJ����\�~�rYѷ:::�J+�b��&s�GQ�g�M�Ǩ�ˣ�Q�3�v�vSu׋���K �����%�T��[�"RBk����9/����zWOC�(�pe$����IM�ޘlbM������A7b����X*F4�B�B�����k#:I�JG3Jy�ӕ�qJt�Wk���-l�b��d�,jͥ����E�]��(��`g�V�u�h*�h��ja�:a_#R�LC����҈p_�AH��~23el���
�\�sn6h�|n�?T�]q]��E��p=
�ŵE����7L؇�̶�M��-�a�M3������������e��\W�^-�����:��5�d�z���j]��T%�Vm�����oo��&uM���9����C��@�BZXiEE��9|__�xNʍ�c ����*;t 	l�'_����#ϐ���с��ʎ��{Z��A��D�^qm�������74fv�v�͝�K^��e�׳Mu%��'}�f�zW�3�*�����Y�KX�=��L ���(��L,-���)��7�1�݈5�������5*^���������?쩏-,���ZI�J�RYU�{��@qV�^v��g8I�>ԩ;�9������[*���~͜�/3N�ժ�|;%&	�G�$%�����co{��� ;��s�|����`�u�C�N黩�DY�a�4fs�s:�i�LG[n#ME0���:�=.}�ڈ!�A�h��Z����H�w�?o��D���rVX�>��.�`�\��meD����u�h���>T+�K�9�v^k/�KtN�<Z��ΎffK�k�YݶQ��T��p�j��)u0ǾV�$�dD�־Q����m��x���������������d��|t�]�����+n��j�˾n��`�gjԺp�>pQi)_ngV��\��@a���»{v6cp}u<������0���_�߹��w���B�*�8��@�q����Z�!�Dnd�������sppE�3M5�pHt����!��@�^f�g�b ������L�
�_,�z���jxqZC0:g�ɋ*3a����U��S�&�z���X����n�òS�P��Y|��W_,���P��܈$CD����<�Z]�� ��b߶[z_�3�K�"p�-TFӺ��u���JwU-$�@��(hGRún��%�8�9 �`��uG�RT����3i�����͌ưp���2���\�$8�`U��l[xggg~������נFTM�{�^��j5/$999�27g9:Hv3	��lD�5������F��+NnVJ���C�5EՔ�py�:fv��Ḇ�Y��s��i����qAT����ƶ^�5R��<~�Ў��2鞃���-c��Y�~��S�}���Z�,���t� R@��aHI���<���nO���"˸7��f�V+=`���I�4�X@��O�����`ᬊ��a���N?{A���������C����}�� �D6]rW�Pa��').T�й2��FQ>Z0݌�C��Q?np%�X��!�+`����dw��Օ�9X���+;��j���!�^/� -��I,U����@l��~2:<\��M�\��Y ���%�*Q�Y�[.:4�w��qQ�q����/�%tb�ɏ��!(=��k�W�\@k6��i� �k�c]�=���՜8��� �3�Gpt�yR��Ү��@n��|�*b����p��z��R�a�A�8I�5�̙�����9D��ӨP��^�05�[�Y��?�it#����L�}�)�I�|~�z�cH�������{1�F��!�=�"(3#�~���B&��Ft־�,8F7,���,
��.���Q1��{���/A���d,4�^���n/�N��>g��6�3�M�[L}T�� ,#��F��s(***�͏<�!�n�|���@��k���(����p��&��XP�ߘ���K-H�h�EC�6���l���/e���~��e֝	����B�L�fͮ�ܨO����L���t�6 �z�]�|L9DZ ��O���M��-C�x;���=ǘ`Ոt�Ȍӷܪ�C��mև@]���L��O=��N�&���S%P ��x�ct����w�ڟ�V�� )殺1������H�q���O��(�K8A�L�
�(�{.׈��F��iC*J31`3�*�/_xY9G3	�6�^�CiF�e�.y�v�k��U`��.�]p����a�ߗ�n��9����ҡ(�����Z���IpK?���u��=lBo�CMMc�n�����=Q�u/��g4��&H{�<�;`�U��cڙ:S8[i��׽H�9,y,q�r:Ur�.m�4�hc;D��.���i4_���h�(.p�)��@+��������W�D}	��ʷ���R�c���h��C/��$d��"�<�����u��g���-��?j��FQύ2��H���%�����l��x�c	�1l����2.h�B��S������RFd����
���1/�����I��1�o���t9����W���]8���,Iud+���Ʊ�����W )�V��W!��٤�D��|?�hG�È\��B^T���p���"d�Rq�&�ݗ��l	Y��z��P�|'��Z�c�{)�����)�Q#�A��d��T͒������>����>���,��ڠ�|x��>�t��9�p�vХi��q��54/���#�js���j�E��[�Sh�S�o�'*�����A��B��~�(G�ňp�d�LA볻�O�Y��h���{u�PL�*���x���$��]��6��TP/7�!C�`V���@�	M=@�`��G�zغx�?��g��L�j���<�h�̧�❗���4���~Q����N.�3��l�.�z�=kD�K9�ì����$���nw�p�M�y�����2~��H0�f'
� (72�+��9ֱ�H��g�� w��|��uO-�U�>�#���<6o��)�f3v�sJ��!l�۳�iw���ǗL���̾����,4SW}rtz�7v��e;���P����n>zd�ª��]<O��'��_��r��>�N6�8��(IU��.�|�n~޻���OaUl�6�&�0�gS��|V+�6W�6��o��]�ĳ���O�˾��pj/��#`_:lˆ߉禖�M���MiD^e��R*<3ݬ�OU���r���VC�U�A���3hD�D���� �>�w��}�=�e���.p��AE{���U7j��S�ވ��':�4zg/F'�_~.P/�+U&t�n彻�"�X�n��|}���vi���*k�u���K0Bv~��Ģ���iD�~n�M��!'�� � Wb��) ��9��Bs��&������U�"7�aeT��f^�n<��u��;Z��y� ��#�'�؉���X]4y?�h.t��6�
�N�`���w8�Ck礼'C����~ק�e4�~T��F�J��F�.��)cP_��>R�/}�����RW�Oq^+�5g��D?�6��et�x�q�`�p	-PӸ���������|ǆ}�.�-T���J��INF�p�ao�g�� ĩEt�(x�V���6���ۋ��D�F622@-�;�J܈��F3�6�X4��������u+Er���)y�Q�JT�|X�hq�e��d�� '���
�a�|L����#��Z��CGe�����w��w��j�)�� Yl(�!B:?H���I�?>��`
�z���O��7'nN�-X@���0a<ν)׬��{F�Ȭ0�vx��»�`o<jx����(1��]T����M��Uu*u��W��!���W'܄^�&i�� ��m�p] �������`9���p�z����l!Y5�#fJ{������!��&P���Tt�'�v�T�]�;F�s0�F��2b�
�f��R>���i&Bi `�=�C��g�B��
���-�q�z? �R��R<5��B��F��	�� ���y�ϜK��s?�ڞS=�J9P�ꆦ�w(�x��3��8�W�Bi@L6���	E��R�E#��
�NН.u,^Q�@��?\O��٠\(�f������ɹ��mQ�����M��'@C���$/����龵Ɠ`��P"˪ B������NEσUA�m-e q��n/�����sщ��肖TH*�`X�Ie��S��˨V��@�.<�H��Ƨ7�'�>�����(�8�h�I.�����?��x X0���⻷ȕO���%����w��"W�y�A�c �5'hc�����f`�c�b Lx�@������/��$��Ye�����u��((b�����J��_�o<"T��9s��¿qt6�R��H6t�2*L4� \D7t���E7�)��Z��X�l��R3/h#�3�����kD&��s\#p����5�5�~�q��]���c�;�Vs�0����w���=�K�Tr���Y~j�-�E��\Lr ϯ�B��d���%sn��;�w� =o��AEÊ��{��lӳ�. e�1ЎZ@�ೠ�.��������!4�m��D�{]7��`r o�,PV���c�4�54��'��rV��0�Iq�h�Ѳj�NG�����'��|��-2Ow�,��+�[Ԛ=_�����-���W0tY�o6�Lwp�Z���h�P<�H�3*E��a{__r�8�*�`ș&gT����h�W���O���nԷ�k�`�Wk��c���pu�D[�e#r�$��'�d��X1"��שTPap�4ތ4�O���v@}�եə!	�Z�S:B'�FA���.c �/JU#lWS{��p���2�~��\���**L��7 \b4G�2Ia)����K=
x��*κ*����U�ڼI���X0p��$��[h�ިZ�p3���8��a�R�.h%f��.����U#�;'K�k�wv6+�Tp,,� �^>]�_,Nc��>�>����.�3���@�T��{�����t��o�啧'��;��"/�3���}��~b����{b��]<�48V_�k�%^�䬚���z��π\h�)6���}�ɗ����f;��n��[��԰p$�eR��h�\	�F��uN�u�i鬚��E%��s(0�B���p ����_7z4�k|_�-�Ч������D��8���U��
��%My]R��i��7��]d��v���5^�����x����%�%jz4�5�kL��m/k�'�ZZ=�݉�	j�;r>��>F
�H?�޲�tTv�f�,��?�w��7��7���?� 1�9X1�8F�^19T��8j���.Lo-��\���J���cP�� �:Z�e[c�Gg���h#0��p�'�t��y���'_���C����+3��t����4�B0�DS/�JE�I�JY�|W���7��r���Nۢ��Rِ���\s
�#_s�B7���b&qkn��K�߷�aV��"Ʌ��G��aS�l%��Ԛ�r�#s/u�P.FGm<�������9�Jٛ�&��fU�c�����P����S���K�s6��Ա������ɗ��f;���{p�?W��~���zݩݑ�tlh���*���Zr�=�7o.�t`'J���KXk8]����5s v�(;u^>�������6�G<�;�����bx��[�gF�O�\5��XZ������ƹx��Ú�D�X]N=3��z"!%EF;��/���\�G��+(���(�C�CD��|D��񣭈��~b_����һ ev���a��o�}98`��Q7\�C�RYS�oOUx�p[\S�޼����~��@�/�
;��XQ�G�%6��wXm]'#�.��@
z>��T�&��,b����c�b��Hw���AG��r~��v>6Ǡ��YblfI��8B����A�M"��)9�Q�`�~��+�ś�|��(%%U��T�c��ڟ��P8��3����_�:GV��Y��?��m�NOUH��?B�+=�rP�F'��34/y����r�ҒQ�r�N���G\

3,k�&�`�H>���fW��Ҁi�'����1�I6MX���͍�ʰD���ϯQ�����v�t�j0�E|��c�|�S�-ۛ�q��]�I%�o9��v>�[8㧴m�a}��k�-S����?��lb�8ρ������P��Z��d:�ۗU���P#�!��x���cJ�Z�S~$�_�[�Iͽ��;8�-"���|њ�hnT�Dhշ,��.K?֧���@w#��E^:�ƝA�]dU��?�[���9�fW�%���Jr^�5��Z��4*�a�7�`�H���P������3��D~L2�7����z� �bwC����X̶Z�+�2��IQ���`����}gvuP�D��!�
t�$���R=�W�iU^!ݒ�Y���.:.&/��N�j�7��C��M�������E�V�p	�@ߦe�&<�8��(�͌��F&�5S}���_&l���ͼ��j|ofe+�:���Xw���Z�dT}����GO!�27b
%=
���N�E6J7/��%/��K���<s�oV���
[�>wv^�O=���K������	�����*kߗ�t�׽1X�L�����všV�S���_��A01�>ѝ4�޳�>������9��3�Ѻ�+�rz�BH,�{W�o~�u�#J�K��/@��W����>�[��o�����cU]O��K��e�3�� ���l
6	����ş_�L�ǐ��|og|�� ��QF��(���8��#)��m>�+�p�n5��'�(�N��)[�J-3( �4
�b�T��O_{57Н"��?�����x���AX�m�y�\�i@��v�p>��Z����Q
9��]x��ːXN��ք��o��>��K���2��z��M��BK�R����vy���uy�����c���7�,`0/����a����dM�>��؞b$�Ӑ��ㆳ!��CS�������|�2�X�N5�ҽ����d��Z��P���3��c�Q���99?Ḟ{�0!�=T]E��sst��0n��\�����3:ݨ������Ƃ�y�B�H�O��(�F��ce�8^)�ļ�p��B��A����	4O�9�cÁ�����A!^-�+�[�m��D���;c�ײ{�q>p,|�ď�����U �����8d�A@~�iޚ��'0>��K�=�^�yT�{�q����1Ғ `aD��%ܓ-�5��\
.gvȮ�2���0��ꪶK;/(��	8��Tnt���Y�N³��\���=wp�q��GO~�YM�wk�t�*��:ʴ5kg�cL��\��t�R;���&�ekw��%%%	�������%�I+)��˧��ptr�S*I>N�n�\P��lO�$���M7hN~��!�^��D5���T�@�Q՘v ?T|�7%㙾CѼ�3�W�0��mg�!=�(z�XIc�O�</�aA��� Vr#F5�`H�4��L�M�%#m�TWW����)�/ӳG	D��ƙs�B}���[#-	P��r���������4�9�f<c�
GF�w��Sr� �>�g�߲tj�q�{ft�89���Jr�����at�n8~�:��N�J&4�0cF�����㹔��p)r^7�(1z��o�H7`����;��WzRD!x�<�+�Iu!��I���~��~�m�O���q�hd͝Dq��!����tH 1���I�n:piG�G4��*�vX1JC�!��	k��Ԡ'�M�_T}>�Va~kg��E��Lf�4Yiy���0Yb~���㓯����ʈ`�w��<�J٩�z�a�le��T�#4�~Ƿ����B���Q���>��E��D������a�8kZ�8E�����n�岹�hL�����A,��Qa��5cYz����*m�$��@�p���I(N��S�;�臎:pLZ���K�X��&����`�w����IL*�9,>`=D�$9X�����EM�<�zM�/u�s���G��R�2=�K~3��*Y����/��A���V�t��5w�)ߊ�ǣ�?e/��� �HqAS�V�F��G:Qa��㒍:�$F��w�d������R���u��x�d���)�g@��-b��_Q����~6�-G�k�\'���ڊ}�Ĕ2������L�Z�,�	��gha���D��VQuŌ���Uv���^wKpj ���Y���g�\S���?79ߵZ�~Bܧ8׈<b5�f���d���P�a����:8���{J�qnB;�\٥�"P�܇��d��8��r:�*���ƺ����Șo��J�pΔ��^���%�n�ǐ�ҟ�NԱ�����){O몁�Q��Os�����0�Wa��(����d�sw��ߏ)
{e�&J�RI�#*��˩Z�}{Y��ׇ�������#�|Vv�<5�O�6	݊c���=߽���Y�N�/$2�˕z����]���i����R0�7l�5:����6�� �p;B������QQ�rƝ%����xB~�Ia�FZ��T�:���Y�7b�����6�m�Ib�qhf�4�o�d� �I��ǁ����;�+��N���p@4�/���z[��e�����I3�`�$��c�Rܳ�V���@��:������8�N�Y[��r����h*�P�8��Wd2����	�W�Ƞy�.���W�y>i���0���??��сl]�?.�B����p������N&)�5�s�3�t�&��[��8y�v�J�����F#���Z�ͼ�k#����`��r
�@��W�8I���ϓ2� ��[|���E?��\E&4��FE/ۙ�-b�#?4"A+��C�K_�͆�k�4��\��S�B�]����(=�Иh�n����C� -�}� (2Ё�z�2R��8n���'|�������@M���Ƀ߱��>}�l6�q���m��z���i*8�wy7>p��()�-�z�iwaɜ�Nh�^��Ya,�O�׺����z�m�x�m��W�Y�mD��_���(`�$�^�4��he\I���$4ysa
���w"$zH�����7� �'����D��6G��:�u;��l��|��l�Z\����Nҵ9���;@^H���6��\����(���R a���`*M� �)%��ٟND�3�9i>���k��Ƞ8�ͽ�[�04�X�WYO�u��szWۋ��Ϯ�|vS���͖�A�3b!������z� E;'`��s:we�Ѣ�<�m9{�����0�a��o�l�{��N�v۳t����3��<5�1e�D�����#:-�r�λW�9c"��a���/�|b3��q���L�aҵ�.�8���p!�$AM!U�����J ;a�nځ?�.E7J�n���	�4~VR��.y@4�ax��R���_��A̙��(�\���7bʄ���ICڶ�τ��<PC(Z��dDg�O�O�X���Ö�8<�Y����WV�.�&�)���m-�-g���v��	���ç����i'�N�e���-���W�r`���D����,����@�)��e���M߿a���$�^�>bM�~��68�XM�ٹ�D�4�vJ��ӯ���c��EZ�o3WPV���۬��Ffep���K���w��m�馫Gs-n�>U#T?�y�-�������5;*��mn��n|�7dfc�I@��]�#��r�;��'��@+�fN�HMA$ԍ5����f8��ѵ�y*;�7�ֲ��}ߣ�/ �)t�#�l�\��L�C���"꯮�r{�/��܂�G�p�RQ����}�}A�B�n���"�)�`T��K;�n~�}"���.�J�p��is���c��AـTX�a�9�eN��D+/��4��wcS��/:_�&ȼ�2��7o�F�Dm#������`��W�k����m���>A������`�~�-T�_��+z����� M��7]�6P���H3x�-�7�~�_}���Őb����tb����)!Hg��=���☟�׌������7�������r�*�@��ɻ�,D����{��`�t��U]�vu�G	Ɉ���۲?r*��<�?�����ct�@D\a��G�}����1��* GԎ$��[ ������ַH���T��9��~���_IDb�j��J���ml�Y>UK槽�t^���ଜc�~ǿ��5:�LP��ǽݿ��[�B���ńV��ן�=}�I��B�3��+���Q-.�mJ�C_�f�=��ʛ����0���B�7��1����:(�(s5���T�OFcM��佻��5�H�t�S|ӆ�F�{̶:h[�!�}�0_��Ekj�[#׮�O2�����1g��l�{���۶�|Y}_tɉPD�4���{tg[8�+j���}��m0�(5�W��D�i�y��0����� �Rdl�C"*o<�͌�i�������@���oh?��n}�٣M��i�iy5E}�} '��k��Y�g�I�����H���,���nO,��he:n��q�	��5ބޏ{�E�k���ɣZ"�x���14����ȉ9|Z\4E���S��'c�;����qAV�d��)��,�C�:�Tf��
~;�����G^�C�[�=6O�^�����E����_�kw+*�b��^��W������wԸ�"������ӲA��<�m� ͎��I�휖�7m9琽�`垵�٭�_���|~��_O�8�N��4֧��L��7Z�*�Ӧ�F݉�F����H�9��;���ޏ���x)�t�=��������X��L�H�����1��V׭Pn4X�&vںO&�;t�ʩ�:B�χ���\+J��ϧtZV�$�3d�}2@M졐�j��9w���o�_�F��X�X����ˇG�Ⴋ��`B�\� �!�s�CL�X���P��弮�/�(�&#�i�_��쏚y��������?�H��{T��/�Y��,{<�\ן��Ͻ�;�gz�u��i��,��< �����%�	z �K�Sل%�B���))i�B�CN>)���JU�\���o�Y��'Lj��7�;�^.�e�}��'�m�LF7y�����uZ�XM���p�s�8�^�������F�����}��'�0dLផ�>͈��n�]�M۳%�����1��Kr9Ƞ􃕋Z��O���
V���I���zD�8��hJ2`<�%>� ��ƴ<6�!�\�F�ls�q�BJ���]��U��ΜX��0�Zo�����(�7nRF�X�6I�r�x�vzOTo�>��:S�T���71��4f��4a�:�,]	��ݲ��
���N�'������l���͍/١&Z=��l��:N	��*:��?�Qj�d5�,~}',�%� �G�%�ħ�`Swm2�k�>:H�z��hqW���[;�eP�㓿��`3��ۗ	Z���߿c��x��zWB����"|������wen����1��5_#"'�(�)\����Gϲ`���N�u(�ܭ���o�,��C��֯�HůnʨrZm���N��YV���^�A�Y���M[BA�=��#�:!47�N�虾���.��&[�����|wA�t(�1<yLa��|�|\Én"�N$��o��Ŝ��C���z�&_�*"�<���Ѭ�W͈e	�����ֻ9}�a��5�,و����
�Y��HL_������1����?5E�|<0:1m���ֹ^US�ȃ�I1�N -4�[}�.>.�X�B��-�E��Fy9�����և�j�$���z� �Tp������?�ݝ�7RT��?8���#�أ�t��\R�Af�ߛ�(7���3j}��/Z5�e9��-�.j���[y�y}<W�Ź9�y�J��x�$���t��h��R��w���g��bB�m���;����'!�/*k�O��Cy�h��֯HzN+�{�"�{4��;�����z��Au���8r���x��[ _�-��}��;�g	��L��u+�����
k"兵�izEe3�Ү>Uy��^���w[��4��i�;N���b����Ѫ��>j���(��A�=]y���s������g�k>ŝ�`r`'�*��K0����Y��MN��%?mk�9�!��K�Vj�ۋ��h:��?6���H�Ώ����M��YŦZ����0V��Y���-^^�&.��G���ƶ�
P���ͩ� L-���.!�r�~��m��*"�'��m\"�؜�����6rx�G�M�~R�>�t�Q�D�t�{�zpdd��qe�V^�q9>?�A�ĩ	��<|�f%V�{�N}��d�00�%ѷ�ۯ��lx&�T���r�����@�����U?\�?���#:)k�i�
>�}�K�Z��c��y���{18��c�_O��ëqV�v�&�۰c�ڂ�(��o2ū�0�t�G÷MJ����Kl��,��KV�λ>K]ύ�_�:P��T��柽�����p��G� s:Ä��%�L�����y��Y�����ь.����h�mK�	�s�q����DAE�_e�hU 0 'O��ߋ�q<���'�u��Ccd��!�u�&�~\�Z����%�w��z���� w?��q�p7�>�d�&6������8TF���x��؆��:�_z0E3X�g�n>�x��<�l��<�"e
7J&�yܴ����g�K��{�BE�l����LlL��l�Z����(,	֛��� 
GBo�ޞn�����h{��њN(.�{���G�d5�-t�*L�l�T0)'��"]��Z��}.&�@v�%���R��~xKvU�|DlZM�-��'JM��S�
����(\����TćwC�Zd�� X��U��#�-��ˏs���^�H��ղ�C�v;B����DBsY{�<>`u��_��gଅ�5��3\��}\H<�X[�������>y��1s���>�w�C&����!��}s��e)���N�x��N>��Yxdw���)��qpdX���$l�=@`13��ɗ�C9_r�����yxCL6�o�&��V�_)r���u0UFd0��)X���i�O�e�;t���~kSf/�p"�	����=NuO8	�m�������)��.�Lxg&�l�ZbTͧ�Ȕ�E#���R�]�ɽ�n?���T��T���]����ȣe�o�P[s{�;������G�	�m'��9﬋����t�X��&Ù]�Cl�u�J�Ư_�L��% ���HC�ih���=ګ;\��QN�'��=��t����㢯�A�w�	��nN����t��m{XߺC<DG�VrH��]���"\���9/�ZF�V^�"{/!�����J�ϲ�9�C뎓��Ob�/�{*o�t��YCoB%� �L��S6��O�TyÝ���ˠ��=־�1�8-�GoX�Oa�)�呯�0M1�N2�9��S��4|���{���G��k�h���<th��G1q��RV������n��L�WU<��3���m������hj��?�j�ܜ��G��1��%���Z��� ���4����A��O��<D|]N�̭n��؇������@��]��F柑��J�(i��d���[�Fo�ϯ�CG��6��u� 	(��d��6��r�2�*�$~���a��E3�����Q���q*w]�,HZ�Kv
�#I��IO�+X��MP��T�w��Q/q���y'{�R{}�ɹ�u��Iw)��Dpf����6��=����XF�L�qm�$�pf���=�m�6Od���WWc���u��v��V�i�"��*|J����S-�sR˜��)ZZ�6:���K�K�4��hM!3���'�)�
��+j�8NI���?��m>]x�QڞaP�#���2 #�4��U�L_��ie��d�QiIC��||o�*;佌�(�N� ���c�E��7���?:����&�n�~	������^��P�Z�����U�Rnf>�Z������+��4�ss�7=����ҥރ�6�a��V�t��a�����tO}	FL�z��T��x�{&�{����i/u�m��N���s��#�p�Ǉ��K5�B���q]�+񸚟�ouX{g2Y8;nT�qt�D-�&�A�iP���ǲ��);bK�bnE��i�D��q��ug!T�g$WUr�j���sV��M�B5�g����ݺρ��m�Y�Y���3e~��&�g*Ř2���1�Xir7�Kf�[w��^կ=���v=�z<\�T'C�H�,s	,���Wa�Y�B�ۚ:r!;ߟ͝�V����+d�U�x�td�\��p�k��v�����و$^B�Ѷ�t�i,�mɆ*�淛LohK?�n_�6�Y8�}v�p��f1E�ch�ٻm�������zIݶn��?�߰d�3���d��K���R�-غ\�Z���W��ʪ�{{
Y��]]�(�o'.Y��v|�C��5#/$���EK<+Z8��j_�b�qn��#��Z	�>Ւy\<X� Frl�L�#\i"���hǌ�3[��$	�,�e�r:~`�����q�T'�A�ii�D�A��l��-�h)��M_oY�P	f:O����x%h��u� �HElQj�%������gSH���˵@p��	��;Ϟ]���5þ)�V���m"�J���a�M�.��Ld��a�ye��Jn�L� ��{W]��� �.�!X�� �����j�"О*��Ț~n���C%�օ�f$�`Tq�Ұ��Y�6�1��H?;fB�����.
�����G���c�&�SD�O}hv㋬)��{;I�u�^Q:��TjX%�ǶlF���5"��"�Z}��[U}�*;D�`+@�sհ���@zb�XVH��+M��r׆�`&XVVO��s<�s(��i��r$�-G�N�a��>�x����"���pd����$*�X��g���mp��#����C��Qq�^x�nF$�,~�����/B�4QaO'��HoM��4l1��
�u���]0�`�����Wr'���k�l�I[ ��\��)|��&�Vt�����
��;�宻������Аp��y*G����0ًIO^֘9>��.���WL6fǽ)���!F8��IQ��v��B�����z3&��R��w����k��x��ď�?��p�2�` ��E�����ſ(�4�q��N�8���|��D��!\Ku-:S�C��ܠ�9\�:�5��@������_�
��0-�G/4>b�VoD���AO��vn��&��1Xts���)�^o��ss ^+�,���up}fDjF�.T�+�٭���k�D͌��%����A�zVB�P ��)�^1@��[&{ǎ����'�$���T6��$�"F�,8��ȃUQ�$�"�A��� X�N��A��3���T��k��0����rH2�}jʖӐ~_���� hB�"V������2�sU	�����˂��%k��ڹ҆&��M��"���E��"h���,bQv,�F��K$Tl]*j5,��=��� ��"H@\��M������Qv�;�l���|���:sf��f��Ήn�7�+g۟%�!@(-a�}�ŀ<x�V,���"D�;�.!�BӤ���7�������^�b�:\�m8ֺt�+{���>�����']'�/O���o�o�(��s\����3,��ڲHr�*뛌_��Ü��jg[�$�$'NìF0�co�t��w!�Z/�dۨ�W�x���P'�o.�^�5���ҏ�UY�d����h�X���s��[�Y�u�O�$,>8�<j��UGe�8ahe�4�������h�[[�3:���j�uM�nd(ݶ�=g��x<���:��YIS�FYj�Jv��xoIܛc2��_��.����̾�F�:H��T��h��������͛7�0�u
�F\ɡ�IA��L���B0�x�ӾE1`�!z:0���}״*p,�1��`\�"����y/hM���o�P%@����8ɯT�-��5�zQJ�j7��(������	;"��eq;��*̙��糒����ޯ��1o���S�tE��d!8�nan��;gd��Z;��պ�T�L�?d�Z��V?7]�B�1����<�2��i�
h�@����i�C�X0�K���Y�o���!=�it��[�d�aogW���&��\���ul��I���ԋ��S�(4�	\�nY$
�J�rl<�ȧ��#)��H8��Q��g���H@��ˆֿ�?�~6 n���������������!���p��
�+&�%�ɗ!� A<�����޿�h�� ���e�4��Z�-�,N��3 6}�����75�3��>ҬQA�'�7���a�?U 7!!�E��>��cB��8��CP�p��%�(���r�ÇrAO�Q���o���4��#��Ę�'ѲTN\���G���J��[˓�3/@�(Cah����8#� U#�\y�P��+L�����������uw�c�M3���5>�.�aYf�z-�Wro���rOqu�
Ғ~n7�R㣞H(Ӑ���,&�#W���V+0��$���X;�\�+**���)̶��mUO\�%��Xw%oZɭ�9al�H<p��{{��c�tь�m�66�7���l.��J�u+Lq��B@
�#iH�T�:ˢǪ�u.��>�:�g���UNm��t��Պ��S�������9���e�e��(�**����P70�����BM�ţ��Ѓ�HG�	�mu���3@>�r��Wr��zՐ�b�䦕�%�KAn��[<�6g����cf]h-��0kj4ffPd�Z��b}�H�*گ$r�,�e��6
3o�����K� 8,mў�R���}~����r��KU��"�UE�@8���ߑ�+��E����Q�Q�>��Zb���PY�)�o����4���q#��.W��,��ܐQ�7�%g���#��6�����P#���^��Yx_���v4���bAyy��3!˘�<�����+qB��b�VWX��Z;�Z��F�Ǫ������Q����(���wl��e�R�o�e �nH(��C(W�|2�l\'�L��e��=k���r]4 ��K�[<�u�l	&7�ĉԶ��v��Q��M��q���T�,_H���Ps��H�͢nU�3�� ���I���n�עE&��P����E��/���<C���{.���t�/�4�F�E5~�H- �Z�RP@�/�߬�x�ր�.���֨�A�8>���ɥ�,�'��c�6�f�����}�θȾ�E�j��W�g<�rp�M���&�}��gd�YZ�n�w�V"�걭M�*ˤ�aQ���p	a9,W!u@���{h�r����sL��݈����|�C��z�7��D���8�;b�I��|Ə
M\���w���a{�
�_��w#�kW�l걣'd��v�� ��az��GC����w#��Z!n�?of�(/�8�"�,�z�"�'��$�A����Gl/��v�ʝ�3��.v���(�I��A��Az��/܈�!!�Z+)+���M�=�i�QY�#��enD y��CU#(�C�֑�2W^�!q���9=Wy�K������:�5���N�y �!�ݾ����)�U
(a�y�����ˇ��'I�4�S���Noep�ʩ�t?Ɯʜ=&m0`h(��?��r5�e]W��������5��&�O*Rb��z�_Lp�^�*��l}+���I�u�z��V���##��O���q�"9ƾ��l>��#i�h�,22��@��L���`)6�c�6g/���;d~�{u��Ç�V�?�����et��n~l�X2��)�%+W{��OX�]���bȹ_؈�1V������w
f��d���f�ʊĺ�g�Z���7�һ���o.i�C��Vu��@
��?8���7Sl�o@������A�-@���G�2'<i;����U޼{����A���ԙB�޼IHv�T�O�6ӑ��9�V���6mg��n���h�z����ӧI�WKC/�T�\:u�y*��&jc���a���Xh�i|�*a.v��	���z�]�X,T��v���l�$�'�ej���(����m���=��`z�"#}�30=�����!�Р���=������������Q�r�@Y!t
]Զ~Å���gL�ϨEi`%�1挃de'�R�8�����xL҅�*{��ut��5e�+�i����'���,91tf�8��-��ѫ-�����)R�P�3���sY�q���dZ�U��e�2>��b�P�Y�U�EIԶB�d����cH����{(���gԆ<���;��?6O��SYiP�~�ۥ����F�h�7� ���٠+�[��X�Agl-�����ݫoUΎ>D]�!�\;�����hiƁ�����{�i�)/���k�Fσ+��y_S浽T�B�:W�W�o�>%9��8<<şlC2��m��;�{Z�{!��vЎ3v�OLp�0�+9�"�Q~�r�{�� O�]bq��"�#Ap�-��Y����|#G�FSQVs�J�� ���M}�L�?���RJ
׵WFRhvȢ##�y]ϟf~�4��_^G��׃�d:���'�����Z���H�sI_����U���ד���tk�5��Umi����\��ʧtqrW���� �Mj6�ѝ{L��}AR&��<Xd�/^�e�|���4�%�����FYn�bY�;;�<��Q���xw��#K�R���ۄd��t5R�'&!6�zU��^�sleclx����;*�"������������C�UUT��<P&��U�($$Td�_�=��vA�K9��h{�X�{��tqH[��z&�d��z����hB~끲b��_��#Z�;�ӉZ�m��eM����By��E+:a툰���!ޱZ�ON�ğ���9�1�vtZ�I�\"i�7#ٕ�A�LBm*`\�8$�9�F�Sŧp}���h�}������z~��ܚbB^�Г`:Ի<�~'�,�a�����@���EQ���ʩ탩S��'l�Id{Z���4s��Ƌ�/�����rz��&0L�2WIO7 O/��v"
|O��)���/4�dzݩ9��~Uo0���[�̼����<Q����Y��^T�No:��Q�ϭ�+rs�o+�����E��+p�.pf/I��L��2�oK��VPH��@��Oi��{mgC!C�Et�}�5�5%H��x;���A�VЃ]�{��m�Z���/I��Њ�k(+J��A�\B�_��hf[4�������M��_|��m�G��|7�)����;f*#I��W�~�������3Pz�j������Y�H��&UC��׸�H���K��n�^���'�&�c�f�ڥ�����M���5����{P�h���|�Q����YV+��%]:�u��`8��_�!��Y�bzx{P��b� 5;融�Ź҂uKWK��菌I�?�(�M��k���O�� R..����
��nx��Fu��]*����{�.�t\���ݻ��y7>�����2�����Թ֞
~?��-�o����ǂ.M[��$HD�Sܼ�t���*lD�NX{�:x+�7`�[J��]W�˦�^�`+q!5�Q2�mM�"b� ����wu�fO^��a��&Ŝ�i�������0�r�sG���I-¤�cR���ÞU�,������ZO��k��Yћnלj� �gk0�A�cq¬��V���J�Rʅ�~���GP����}u)��{��?���>�Q5�^T[���W�M�;�oӧ��Զ�����������Ϸ���;p�/YZ��R����:�����jv9Nwi�2,|����$�k��"�۲��3n����o*�x���n�/�r3�Ԧ�IP�-�ީ�dUgQۂ�fی��"X������NA%_��Oϥ=���A�������{��
Xⰶ�Z�c˹r��������[�]��4Gʕ�������ή��¬��!t7YK$&��T+U~���u�$H)�^t�$~W��O�S�c,^x�~���{9����/��S/������7���V/�O[�����7�oPߠ�A}�������|���)��S��O|ۉe�!;.�p�<�M��W�)�͕���W6U�z�=��`�7a6dnyPf���f����y��PK   �n'Y���n� 6 /   images/ebd5c09d-583c-48f4-aaf0-071f49184249.png�eWA�-�܂�ww��Ipw	�KH���]���2���.���`o�u��<��p>���kU�޽�v_W�U�_��1PIP߽{��� �������\Ȉ�"�{?k�5�=4��UO��{�面����ɟί��˾�M^�����.�<DER��	*�3pƞ��щri������cM��sE���F��xvѼ$q>I~C�����s��Һ;b��x�.!aRn�xa�~����[v�D�3ǮEփg�#x�SG��d%R+�Cm�õ�!����^�q��|�:�ڞ��/�Y�Q/X�������T�|�?w���Yg(hZ�l�o�������o��7�Kx(����Rn����/�v����J>�Q#'���?J���D��+fV���Ob)ۃs���!�鿬��� ��.�k�?Jb ׳��a�O��o�O��'����W"t�aMxu��C1��|�5���@�N\�N���C��9��veY,�KR�s���QϷC����ofZ�E�������z���禈e�7��;B!B��䘑P�aB�h�H�o3�G�ʭ=\��4�o;I+pY�i\��(�!���9?u��,BSC@�:8������Xx���`ܟ�l��'�WE�4�U5�W�ur��*h9X`>�:D`g��yR�ǖ�_��iQ:��e��Sl�A����V���Dz�l/�9"�{��K���X��[5 �9�$Ut�t���`�h�ۥ؎�^RG2`��С�|�����s��@Y?�&��M$����rt�棸��F�K/��ճ+fV��Dk���`p5�NDs5G��fi(|~�Y�<��:P	��lv�2l�G^_�Yy��������`��
V�j��ؼ��E.h�ZJ�4bH)�fh�c�&��j��FS)���O�7�|��T�N��6g+��jX���~��;K���1X���5LL�}��1��,"��n4{?��\�KEp�l+�l���;�J�$XgUՅ̹u��sN%�P��,��k�!���l��:/&a"��}I6H��$e���J�"K�b!�wz����0eV%��K�y2J�)(�h���oZs�u�%@M`�np�ܙڋ�=����2���G_��.��R�>|��&&gR���� "J��+wW�����ɱ��+=Z�<���k9�ϻ�K�rq�-_b��!Dd�[��F����%!,B��_�6�'��=�b���mI�^9Ƹ������R�LX�p2'�ٙ�qy�-��v��?vI����t�#	֦Vc��Ո�s���J7��]�H$���B;�a���j�1y������iי���F�l�y�;�ԏ�J�jpM�](M��@�u;����4��]��	D�[p���S(B2,�1��Y��iZ�ob�u �U[ŕ��$��s����<��cP��gr$�+���fBG�hj� �:���tt��}��ƆYހB�ม�׷(����U���R���x�Zuq���?fbCI�����*�^�Y!����^��Vk��S���<���7w1[���:$�m%�d��X�Z(Nھۓ�J�l��F�QH?�lt����V� �2�����_�*L����,.���ݫ.�_�>��E�l4�����[�1�~�{��wjA  �E�4
0T��'q���DjT�����xF(��E�h��I7��2�8v��7!/v^E�+<�M�{*H��8��DRRr���5p�g��e�5�pFUBwI$S��%8|����S �*�gx��)�= ����2R[5߾���l��g��H*c�X�2�A�U�YY'V�_�S,"��Q�K2�T9%΁�iϵ����koêOgq�KWk:��'���J(� �S&�����$9eR�6L��Ɯ8��A��&��?gN�D.繨~I��D�L��j�p�O_t͹�6o��,�����xտJI����WƐ����*�z�]�"	'�ja�0�Z>�uY���N}	�`D��g��u�A;�@�}��{����c��gi+(?(�^R����9vxIb'���9���=�Q�j:�w�x�&�m'��W6�u�X��˧cvkY��l���˳,
���"M�Bg}���Fe�F�N;*��r�m�0ݑ�2:X�����A=��h��Z�?
@Ér�$E�a�v�?e-I�~�&������KrE`�/��Y m���������0���Y�����`��p<��8uͬ��\?"�OV�.�r�:��� ��0���z�ܰn���̯���x2p�4n��ߨW{�C6���`5���q��O��62q[;S�lfx�ʇ����HR�ك[z��h�J#˔�\'T�m��_8��̓������<��rG|Z;!�Ng$�&v�Ce-A��w�.�[#Fǀ��Т	�j
J�����Rݙ��E��eg��;q��v��u*���Bg�#x:�n���TM�g��h������0Z)�,6�2��w���?׼
���zZ�C3=����3p�(��U��j���2�
X�NQ��X��&3Yy�3���Kv�C���3y��/g"`��t���[<����DW,�D�4IQ����.��4���}/TW��sk�~��]�7<G6����՘�ap-^7?��n�DE�Qu�n<���6�s�gF�=_��_N]@5�7?�v�#�1w�HD����n�wp��.���������k*���ϙ�0���(~�BL�`����j4;�<���Bj�v�q�=3��x�^v˒Q�v�\g��A{s~|�j�f�ܱV��~�U�H"K'UA�JP�8d��4#CP��7��7��7>54� }�,��%g��AZ�˦�룡)�k�����ꖿwb}��*&�=�3IJbN���`� �X9�mv��O����pvt��ZJ�h�!�s��6A�x�qw�А���>���=����5}�QXl��¨UQ�`5v��]�uUɏqXzw���c��=���~�ˏ���z���:����Sb�ʔp��N��bK�����~�P�(�u+�*aƨQ,�$8���0dD��q3��Ȥ�rl4^Ř <����f���#1�|�"ǅ��ut�ajN�f�D�Hur�',���L���	��
^��Oq�����q��cV�M����_ڇkT	|R� ��&�����c�%��D(C\����YKX��ZY+�ܶ�[�$%�L�L�G ��WO^?�p:D�%�}H���|ڮp�'���QZcѭ�Y����Þ�����%՞����/����8���3sl�\�d�_{7N�M���\����8�9�/���Ī�}��z� U0����4WWo��>
��l���^HFG���Z	{G"��QWpW0[�M� �6s�Th�s^H-&�Ì������)�������9RS���~���Y�%����h���*V�7���e!Vv�#�M�� ��m|t������4,q���V�k	
��8mLTB	Z�;I�;7B)�f$�De����{ǜf�d*��(:o} Z7��.a�n�埶��ph�z�j�;���H�y��0��/�813�l� zͱ�O��s�<�l�?Rk��4��"a�[��}�S��x0�U�8�YVVWg�F�i�D�����U�Jj�IC�����o��r���߷��9{��0��B���\�Q�
i+If�{�8/��27�G-�2;�ζ[E�O�$���R��,u˟�~��A��ݻ��%�z���S����-Q��ݥSԷ.����M?�qRs�I`{&�;��5o|6�ǿ�T���˯�
�)�ލ��/�*B�`����2����O�'[����=�}���'�e�9!a��P��*�y~�|4_���<�r)�t��aP�QǗ=@��ۡ�/>b@q��T�Z�\I���ڢ��e��W�����hw5�hneM&�)CzC�\*^�����}2��I�Vsh4����h�q$&6�-��%%� �����IX��cb�$�y��ݺ� ���
q�%`�:S� ~��IJ�DF:&rH�@�;'�*ƈ>�)	O�m4��,"]��O�4§�<�R���^����)��ԢJBr̻gx���m�a�X�v� �)i�:׶��,�V�]�¹RlLh�V�K�ѽ���;d�3g!���{�ҩ��vBX�[�G���uy
_��՛��'l9�����1�8'��T@���|=�t�p�W��T��O�WC��#�ſ�k����_8�Z�k�l;��ᦻǱ!�I	�,W�2�!�"��r��ӕ�?�H�8�Va���W���5��ߒ�����]�G����UA���h��qg����Ѭ�Ӌ�����eMl�,�N(�V�(^����D_N�3��Z5}���O�}לM�b�>䞊5\�.Ŋ�)�e��HT�,^��)��<-'1� [<���T�Kw��!J��#��q<#h*_yૐi9����8�{ɂl��׷�̓��-dW|��?½t
5ơ��H�[j&�"��Ĕ�E%� -l��h�M�o���<���FGU����&��ڏ�G *x:kEL��V�q�-DIp+�?�뤥��C�Tf��P�d�7R�V3�1OS�$���V�v��إ��]Ss�����F	����ΰ����a�����þ�d�Fkb���M�TiՂncE��c��ݫist�����&G5'���G҄(-�����I?��w�l]țs��&��.Q����p�eА�����7�x�Q�F����6�wv\���h��
J�����6��xY�=��
����Aa[E�u;Zoe��O5����5�b6�'�!�a�յ�5V�� ��R�|f,�] $�ăZ�� u8kԑq؀Vc��
��G���Zˁ
��s����G ����� rmk��ϣ��m�(S;a�*�"����u�_���,�)�f�l3d3��9��&-ݿR�͜4�J�D*�����2L�щ$+ t|o�'<gc�)8���:uB���Z�t D�mKz�|#��j�ǝ"�"p�G��mq~�J�?�p�������hly���r��pQ�!�b�m���݋����吋p�~5�^�<���D�����X�?�}(���ٷo�(�ec�t���찭F��Bur����S$ߣg��R[zU>���{�\��g��7VK���A�+�g�h����k�Ma��/3J�2F>���/�N�r���ʿgFEMm(�����☘`r�%�_l�8s*����j�Q���2,�'`������]�+(g`E~1^<��d-�1������
�b���u�@����\/�������Za��P�3�KYF���4k�KQ ����wF�X�k>j�]*!�呎�k��9�(�AO%`4�e�4jSD��"��3ӎ�`PK/b��Ya�8Ї�uv�V@k�g��wEYT���p��x����[_�(����${�k>g��+.Ըk:8�{pjA8(���Y1��J�pR%�H���?����i�Z}������?�f�|c�VTu�������.8w}�s`�ކ�[U�
;Jy���ol{X}{�*�}����6���LJ�}�7��y#����yf<e��iw�j��8d��S��ٴ+���^s{iɠMڢk�o��/�[���0a��Ta�����'�;�X�\���A�[`�(Q��9ZP�<2Q�mz�[&���.���;�Ζ$�B�Z��mڌhʒv�h���U���\��r�:�j̮�^R�)�W_\����T�v�my�cާ�Y���N�q;�-<�~N��� �Ze5張>�K�G���|��\ʌ�~���_eJ֫��e��;o�����@Sw�}=������a�ZJb-�b�EAri)Zee��٦���:ŝn#R`Һ�$�T�Z�o��O�OV��>2�(n���6H������ٶE����o{Rit�F`���3/&u���r���C����L�T���mCh�AJ�aj(��g1Bv't���Y�N�F��]��je�^=c�l�[��Z��6g�!y-��*@�:�/-̣�[���i�e���� h#�9��x�g�9�����0e�f�r���)�2�+Ry3&� �>����B�:�z���v�""��c�B�9�j[��ė��7JL}ޞ6��>|���:����	��'��:�Y��T{BF{���ٞz�!�����k-֎)��T`!|g3���Ԥ�n���z�Gb�~/s%���n�i�.i����.���7�Q��B���'g_%cS��h) ����QDSo{,�Ö��z��<���0�!	�� V&gJ���Z�)�c��j�~����]�8�dNT���9Wڙk7�m6M"���T>=7����mcBq��l�g�Wl����\�_�%GR��V��>�Q������yQrS��/�j$⒗R1 6�Z�'{{�V����L��-ĺ�+�2���H�ؠ�g�Cp�Oi�H�4v[�h�ƿܚ���h�����7���L�4ݝ����=[m� ���4y��Ǣёbw�q{�m�x���(h��H�US�ڊl[����0�:P���Sl"	����3|s	=�Jr	7P�r"�{����i�&|dM-L��p���Ն����!v�m[�b���XZ��S1�ƺ�ď���-��O�N�;��t�0 �O�����_q�y��|�p=A?d7Sǿ(pmUd�g��P]���
ʧA�\���_�Ɛ%������w!�D"�2��	��T8��[Bi�Uڿ�N9���]ՙ:��O���e^�h.�2�.�����W�j���U>��	�#�<2�vo緃��0��W�{�����z�T�����c2p��gV<W���B�-Y{�-\{�~�7>Lz�+��1�>2�F��f�0�ڤ���r�}ܼ�?���Y:��� Dz���biP+-�������0M�t/Ag��a��^��v�>��y�r��k�<]o.<��?I;@Z��|�q��镖�=+Ǌ�����i��q����%�"�-��N�1>��ǳ�$X�Tf�ݲ˔����$]�rE���U����$�L��Y07l���SY�Y�@m�US�(m*[-k��%/����\<�w.�fA���Y�,b�M��
=;坈.`�)�?��2���(}m��>S#��Tx�|̝��r�T��y*��'5��W���,ۃ3;�K�4E6'%3�򱖖/�;=O����Z:8�ψ�ߌ�)�y%�h��1�����k����R�xK�uo�U?�X���, ��c��_���.jB�/5�*�����������Zz���B��"d��I��sL[��� ��?t��(E�U�u�YujK��w�[���	���z�ְsQ��-4&=JAd����U�n�p�X�q�L���@I`�b�(?!����Z!��H"3�@$�[���k��p��Y��#�0K;)�w&�씣���ڢ6�1��dL��> ���>&�+VqV1;�YĐ����K�����Uf��f��h�Y�\�"e,mn83��+>-�<G�+�oڭ���r�޺�%��Rb�����6$���x��q�����������/U"�P�����:a����dߙEྷ�1���{{Si�I:oZ�=�M������Gٷ��G:%� ��p����b�g~�O$�G���W�r���CB,�h\��C��E�iF�Zx���s$Rh'�����RdSb]3�m#�Tȹ^�.�5�����/�Rc���-[)-O�͙(@�["-��};~��і�)oÀO/g����D� /�L���I��:�z,�*�2'����w=�2�+��>��~9��ر?��P�mw�22[���R�:��Ň&�?���qޛK:��R�Tn��C�Y��YL�\���C��UJ�8���I�0tT�?�s�^�f��j�-���iY��V���Z�0g�*�~>�=�� ݕ�՝9�C��V�t�U����P����$yơ4��P6Z�A��6�ݭu%GZi�]�l��ڡA�le_?�r+��(�e��G�����*ȾJ����8�@]����x�l�|^�,��4�%����9�Ūr��p����jH��i�|��S����1|����Eə�����/��爲���[xL;� _	���1��f��R	���E�egL[�pr�%zE'@�׍�);�_�|�I����~�[�Z��@������r�O�p�|�Z����_��|yW����}/\�xr���5��>�#S%њ��X I�۬"�bp]K�WʘOWd��=��y�H :�EK���)na�o��F�f*�%I;��*���X1l�GI�Z�z��3�:��T�\��7k�3������|r�VM��@A�f �"@�����+ӎ5�A��g��'� �ɒ6Q�����mǏ���mm�&��r�b�s["�UV��a��́@�Յ{�v/��?(|�?���a�a�p��a�7�����A֕�-GoP�.vB��_�%�'#�5�o�j���8�׹��0}e�>V-�ݨ���>��]P�X���2��|2�&�;��Y�M츬F����2�_�Sܾ�ȷ�[�]]v�r��w�|k!?���.�ʗ�W��E6�C����Đ��'+]G�ൕ:.���9ɻ~�5;��U4L�(*� A�I���&������:F���F^?%pCtclUg㘴Z���D� �X�s�_k���e��e!ȉ�|b��?�6*�F��e���;�ַuL�#a3��y����#���*��P&�������Gk*��"�c���B^�
K���c<�Z9�?8/Ds���Z���~��/m��~�ES�D OK4G��N�%v�����O��"i�����IQ�X[���� �Мxź�'V�|f���P��\q��P�>M�����	[���8��Tz5Ǡ&>�� �wz9i�P�ӟF�����<i<ٺz�fR#�!�ȯ������ݯ��ٵ���u�]:w>`[Q�k1���+�����ޮH��������(�N�E6*���,#���1��ޢ¿]d�����%L��o�f��c�_��K���J,�_�;g�`���W�M�Kk�u5�v��I�3f񣣦���.��;�
8��+�?���w�${mb�p�Hnw	���A���I⡷�.#P��� ~P<V�چ��+ļ��pQAo�_p�(uTbpfn%z�i��͕o8X{wi��t!=�U�T�4�{-.��T78��T3<��.a�PA�<�-q��V�R�������ՒF;N���u
5�+����˚K���j�s�ڮ������e��ֳB/�G�#�9���mg)㠥�Ӆ������bn0�A���e��Wf��#l�VN3� ,��)Gn+�~ՙ.n+�EOe/��������[�Lsm��i��"/�U
��@���A-Z�Y�r��Q�X(|��!Y'ev�B{� h�J����|*WL�X�!�q�?&e����#$�0�G�#5O��������r��)���vs�������	Y�V\F�d��>�xp$��	���Dc)���AY�/G!�P��]�;�$�c0n>�>�X��G���n���
�^�e��y:
��D��Xڍ�@�J�4���;�΍ѹ����z�3��B��xA��I�:`��˟���!o���	�O�J�Z������?��A��}��٧b��S��}� ��О0�.W�����G F�KvƯR����}�Vn���$�ĺ^øx7�6��'��23��R����qb����� M�2��u�����]�B�(&����@����qOlU�7`M�k:�L��PdH�e���k	�G[�uv��)ko@h�����2����r1I.Qݴ�&� ���Q;0_��m&�����j��Ѵ�ZA�o�g� �O�WQ����=���"4��<�B���bp�.c�x�� h�У�;<�"Q�674hfw��~�C
z���w���{z���w9��=�z����1����2P��
n�O����( �}�-�;���Dk�N��֕K�NXT*Q�lЇ/+qP������?��r�i�<%��l����ʓ�E�|v?���J�{|l��VqC����p��=��q{�����y�w����	$�=�8ѻ2����ј����S&=������o�,�c��ǧ)�����l}㏏�%m���I3�h�D�(-	�q�Z#�����LZ1�r�*�Ӯ��։�*i]�;�1;�����6�� �のs:3-�%>�i�v>�6!H�;;�A��q8�����O��đ1��><��.��LX�������O\N�:��S�)��4���<lt,ŷL&�I�_7��*N��V�k��.5��f�� �V%�g���䰙�4P\�o+�AX�ޯ�f��.u_=R�˝�o��Nn���Ͽ��yp���k!�
�2N/�s_���u�mPO�h$}��yUo:��7}���.[�F�P��ѡ�SYQ�>�B.��(a�Os�-�m#�����Ǯ�\���8�|�a��TvApS���M���ho�Kݱ(�L�o��ON^.=f��qÈJ��y<C}cfŐ�m�tg�2[��)�(9X}G(���.�p���]��jt�*�ʴ8VR,��J�#p�^����R�v�:�am�욖�>Z+OYQ~�Jh(�Rol��ш���ę���0��#D������;�4�=�2y�D�����/M���cŒ�#쳀P(����lv�D�/�^���>G0D~2�d��Y�gL̾cO�\�D����ӟ$�S�ti�	[�"=�{�뒕��:���
���] p{'���K���m&T�jOw�\�a���)���s���m�k%�\��V�\p(�;ɍ�vs�W�:x��fԀK��^.���oW1�B$`A�A���m�w6�"���S�67���<I݌��1������Hs-���
�v`M0z�X0�-����$D��R��Q)G'�Y!W���C�w�G(�ȉ�tR�o3�Z_�g�'�m�;�)����7���`�]ߐ��W	5cя�Ó�S*����3�}�������|�!����M�چ�IՀU4*#?5�������0�b�6���UA� ���P,m}-|���!��0��D���G����DZE�����y��292`�GvA9I�j�^X����G�{ES|`9�@Y�=/�E����,�l��W��ìw����G����!�zl�a�7���0���z���ʙ+=X�B,C(f�^#M)��luj[��n��u�.x�ՠ�[R�m�e)��!���Ѡ��p�x�����i�g�@t���L��~�ᴓ��S�Y�/LӴK7[�D�'0��S��.�+�㉮����Ϯ�гr�D�[�E6h��n���͛>֍K�������ҡ��ρ� //	N��S��U .M���n����俙8�$�L������?�H���3('s�2���~��.͏�����d`��\��-I��ͨ�����X�' ���,a�W�RGa���ի���$�)�my�X��
��uU&�����g���������rf�J�#�ggWz�5%�/���i֨󑑸�Ll���i}�F 7�$��9�������
��3�4.r�M�ȹ��q;	"����</(S����Np�\����=Yu�F��C:�zt��o�V/'j�Lo#�a�U��L���x�u?�]�v9�-N����y��^R�_�_�E��6����u���]�k ����;gr�Zs�%K�ʸ޷�3u��G��;�d5ْ6�솿�sB&�Z�[>�k�_�d�+��/��C��]��
z�J\�B-i�������T�o���%��"Znd$�_�
~�������Lw�3��:���[�^]e�e�2p,�r�>�ݏm�ܠcz��o����Q����1'�).�(���l>�׮��~B��q�~ ���7	b��3�ſ4�̱�ƍJ��2im���(�U�A��fyb/�w��H,���z��ȪӅD��p<<�^��]m5�ٝ�<L��	�iEK�?Q�f ���N�&�\ұ0�_��5��U|'��'����v3��*PT�9J-ӄ)�VS����y�8�u��і9T�M7�Y��`�����(�C��5��f@Lm����7)��<��Q���w҉���'끢�% ftĭZ���:u��(A�mm���*��հ������g�)��u�M��<ڎ:R�D��j��Z'��;����w:�rd��ck�n
Uq�ީM��b�/����5`�I��u�v`��{���U��Ü������sJ���s��ٌr,Cs����m�T@�Ax��J�@(+@Q;����A����e�q��"v�ZNf�~܊i����\~�C��$���A]�6��NI�Ka�Yl"6+�(_˫A���(4��Rlc}%ܒ��G����H��^�B� �ܥ�W��٢[���v����s�Bj�Z�\�4V8��N
���>���$�
��0�2���-���v��D��ph/�s����J���7�{ݏ�v��{(��و��E��Tu����U�j���`#������h�h��7>A����d嵥M�,4���[:� �zv�v��y&O��v��}����ҽ��� �t$������IM�~�EOៅ8��u.�O�RZ1'Q��@�
%���:���" 8����6���W�`^2�H!�Y��E�Sˤ1]E�g�As���Lv�z�W��O��X,4�`����~G�����z��Φ�|�
3J���o
�"�C<����+�s�w�}�&�k�.-� W���t�f�P$l��s�����e���1���Ie<�G��yD(O������VV�Sʱ/�J�����������\Nx��?S��ޭ�uZ���rk9=�GŇ�D�WX�$3Ԧ3Џ��%Y	�%55t��M�߄`fz7J�{=ћJr��h?���|�-6Q�ξ/},��G�JYf����p�`�k1ӛ]�3�|7:�z���xHp�jm�*��0`E�RЃ]S���*��������7z�f=>,�Ѡ�z��ܭ���c����v`&{�f�@�\6��S�A#w�PGdV�p�2��S���`1���g	S�X�C6(@^_GB�o	4nV�o�)���Lp����zǘ=��i��-���՞�vL�3"�~���N�(ȯ��UEq�X�SIx,���O>*�;�o%��aϾ��*6��qH\�
2��������SK
AÓg�N��m�/��>���<�s%����L�i0Cߥ �����By�샒�dV�|�.ض�13��C�&� m� P��4�4;����9#՗�3�aL��q��į��X�)PmJ�d)�>/]O��D
�C�b��Q���[R�i����4����H� �^��=�_�'�oR�t<>�v�Pn�wDU����X������)y�Gb3^���� ����o�WlØy5��L�nې^t�mj����'V���/�nO�/���ɰ4� �P�u��u���|��v����M�g8�cB��W��4bDP�<�J���+��.�����cF^皩��nuџ___~��$14"�a>�P�ru�,,��v���X�e�3Wy�������!߷f]B�i��*Akp�6ZQ�'p�7M=X��c���+�i	ڧ�p������h|E��Ssxʹ��E1�drO�����ܙ������Ѣ�\������E�۶� e�ݜ�*�	��K锹%g�gpT8J�l������B�]R�����gRJ��i�ߎ-˴�l���TVK<uA�B�>����X)B+�!_w�o�׃����m�}r������>�*��$�l���=y��� �����yf������V��w3,J�.�*�'V����ucC�٣uR].}D��UܞTQ�Lz�w���Cmﾟ������J/�s=z
�~R�̯+%�؍B5c���H���ׁ�X�#��Vs�������V���L+[4(n�u�3N	�F�����!G��	��@.�����N���)��Y�->c`x�A�O;�XVY����{�[Q5����j�>�~�J�z�Pe�Ɠ4x�b͒�ah)�s�{̢��p���Ρ5��pr����V�R�g��"�kffJ��Y�E���#k�}�ؼ4��ϳ5���!�b�nf噲يS�E�T_
��'EQ�#	wX,���C[��I������l_ǁ����
��H_�Ry�|]1�k��yK��D�\w
25�?���Q�1m���t�gyY����@N��\�qQ�3��r�#�#�"�����>��̇�̑��я�[���pL���Ρ��"I�l���Z��(��t���S:Fީ�ʘհ�Us#V��R-&"51 K��;�Ͳ�I�E�c�H�I9lu7n�����Em�q�m���W��nt�11�M�L8L��XM�����1��Î�v����7��5	H�]U�=C�.?��֚����8�ⴷ��K��$r��ye��EPt��u�Um�@#��z铐���h�s	�z/q��2X�\1e��v��\��H/f���ښ���/�3��}:�g�p�w#xT�o�vd��Ψ���PG*O�l���`��b?==�ٯd�w�� {�J�mIK� m��l�RD����F������n؆*b��˛ƾ��1���>Lk�o��e˧$�c߆���=�<�go �L��K#�O򷫗��#i�R�ٷ<U{��?y������@��3��A�&������U=�׈�����Ƽ�����g��?#}�&8���{ا8.n�[�k&n��s�yDa$��EW���s� U��c$ �gWX�:U��B�wbz��Z���e$�	QM���⒊���֪��x}����H�J��՝�&b;\jl�'ޒ��e�p%0=+6��6�,��`�yk�
aݶ�Sg�����/=��]i�q�in8H����sQՈ	�ś(�r�,����D���f�<,��I�/�҉z��^;t��ϞքTvg=]+� ��8��@��S�ρ|��g�߂��]���k��QG��5<�u��ɕ��7���ɛ�GHZ�z�z*��~��8E�nz�KU	���N�}��Ң�"���H�^_���I�w��j�g�M4��T��jK�O��4����X�t+;�ғ��2�&ԕ�պ\_����}l�����5]�щuf��D�g�3���d��;���:
;29�uFd$����x��#井���ͼ-��I��:�i�4#�Ɍ�+va����� ��g�0��^�$�0�[�b���3!d���2�ߜ�{ R�������G�b���P���?��#�ZFy��tџֶ~7aR#���ԫ$ ��^"x?U�{S���Y�8`��I��]
�۠G�s���M�u��ӦX� b�^F�3�K B@�N�l+D��tʴ�G��g����G�`�>PA�;���h���D��7mCWD2��=8P"%�̣g�4�"�}�cr�"�l���n� �>G\�2���U*5��WG�m�+.�AF]�O�zO�Q�E����Q���K�s��?�.��:�%^P�l��)Dz��:|3{�>���:m���{#�vrɟ��nHn	F9&��Ks�0w����n��?�t�����/�'&��IR^tĦ����P� O�AV�ً����b5�@�>W�˾0p$�S9E�OS�%��f���'��RP"��P��md��r�0�dwz��^����NG��ɱO�5g�p��\/��qNn�e0^N;���i�@.�zׂ>����R�k�gD5��n�i��
"��[� ���͂U�ܶ���L�,�[7w�[��ȅ����C������\fn�l���1��"��
[g!#�\����.�.�������<��I�[5(�A-~�sR��(�ƮpSM�����z��/F�7����X�z%8����,!�O�� ��֍�P���S<�:G{���>��'��fyG��M�/��c�c�-9d�֘z��:��C&~/�S�cϵ�ӗ��O���Ie5��vKz�Ը6�#��@q�����Wzb��5�5}�>I#c�͞�2^��&
_���A%��%a?	��4��ݲ��G-wq���eM�x
���y��=�!b���k��H/~�:]��Q���x�"`^'��06}+bwӿ%����Q���`�D���&4���c?�ݴa������$SI�=�*���x���js�%�j,�e^f>������������߰���`��lWzue�zi�G(t����#�f�i�Po�8�
6�!z��������zЙ% �ɝ����iy�`x1���e��	e/�� (@׿��41�Sg����.���������Ȕ-���»��6�[&;f^����C�	?@75<T8�1�ɓ'M��oݽ������s!�EK��&�
��<�{;h(�p��4�UYb\���+h51������\����?���?��V��l���W7P����S���<���a������F����A�A{��I���}��ӿ���ĳ��O?��EH*J�[�+��GQSmͭ�' �-�HVzNIb�	�����'���4y�(Fkփec��e��DOcKw��l��N�'i�ԡ>L�4ej��U�D,r����i��Z<*�����ݗt^�f����{�B7d��zA���)ǣ0ݯ��U�����,YJ����s
u��/�%�������Dm�6���	A�3��O����Ԍ1[�^��qcsm��M�@h�������!���l�i�5�*���S����"�u�'B3O�?�	�mg]'���>�t�w�7fNH  �B)�@L!
���J���%T-�\�vWk�t�����]ݖ.KJ��HBf2��7w��<�����{�wr}I$��ﬕ�w�=����?���[0������S�_����usS-��Q	�H��h�_���(x������eg���CM��������g�!����?=��=�sQ$��
��zQ%��Pu�./���� ����ޯ�Ӎ\]QJo�R1/mWn��Dc&�XN6��.J�DI�a�jZg��"�PCV_m�.bb���M1z�w��PZ<�,	�2u����	-f�����p�3
jI��MG��Is�<T^O� !?ub�%0���j�.��KeD�x�H�a|��Qk�R!�=��+�Kޑ��玢�7M3p]7�?��:�1�C����N�;�B��q�Q�oEaܜ��������l��Cw��p��|x�]w5���s>D���?��c_��ǚ�N��Vf5���U��+P�܄��!<�1�oL!W���"o��zIb��Z��3��ôm9Ģ�ž�
yK㐟���`LDw1�Z�ڜ�u%yJڂT��!ș�Kn�p��z�S����� �%�K/I�يu]��Oň�jl�6�q����|'�x�8yߗ�r�q���S�+�a�f��xj}|���<��ڐdm~jJ�p�����:CF����O�ѥ.���9�sW!�r�T�5�~7V᫶�3DD� �B�;2�M�3��@�2�7i��f�c�m��u&�L>9� �V��濳Y7�$�2�[��p��CL�]��, g����(�${W�ƊT�L��� �cI�}I�p�
CIR�ቼH�4�	5��J!�����h$I7y�Pts���X\����� K���!���|o�d,����4=�U�s�Ц�&R��g��(!�>�H�3E���3�������^�3rۦ��)8������ó����h�Ch+Á�����7{A��0��������O�I���PY���r�N���|��3=c;y�,+��i[8{L�F$�e�D��
�i�U���(	�k8~�=ݣ�esZQ͢7֨~� Y��S)A.ެB��T��\�ʢ�J�O�l�2#�(:_+�BZC~��i �� ��}ٔl����"��#�q6D��x>[W��>U�X%�l����&[�q� L毒��B!��z�rˆ����mc�K@N ��7�i��B./-"�/�]ڻ<�x�l\O�\'j��a�*�q��i�N��3����0��k�J��(������0B�ʝ�T��nj�ƨ����\n�X.SQ��L�����޿o�+s�|�{N�w߇׹���mE�i��fe�i���P��h�|�g�D>����ǥ}w��8s�<�|*�pTs)�Q����h唤��%�FZN>���C�� ���P\"��:vG��-C�;+XEq�>hI𕖪P� ;u�#�x���w0g��~?��eG���#8�ȃ�}��C��Eiz
��T����ŨXĉ�-t�}\�G�T�S�63W(�X��?�q\��w����ë��%�����>y�U�P�bݒ@�)to(�j�2o���\O/�9_M�B��P��čJl�SA��9��h��ئ�'���~V����t:\Kƚ���S���@~���������F�" �K�*��%�����3�'���p�}LW�p;ۈ�D�	 )~���	Vtƒ�˹��Q���̱+oa$ V�@�&�En=�0�S�GD2ڡ3g¬d�N$$O�]9�-obC��}X�VR~S	aSJ�t�^�o��N�\x�d��}�+n}�5�����oto�]���|���W�=�A�~�e�sY[33��K�"�lgԊ�Z�lŲ*PZ,2/M�O�I<y]�x�&�8��d��?'�s����|6� ���R�i�I����B����yN��C��3����pk�8���Ya�;Je�m<��/V}�@#��F"��XG@i'4p�JW�M���v`X9�Ʈ��I����4;:ɰ5�$�I�*39�]�f"�U9��
�r���)P�D\2 ��� �x��*b f��À^��|)u�I��r��~��t�A	��oR��]�q@q %]�}���Tq����Ҭ���;���ٹ-˲��e_(�
�r�ܬ5J�Z�թ�Y�T8=mǹ\��\2���y����{�ڃ޵z��?][Z�[:�,La5?�N�
��xZ�Y��?C�Iwr�p�v��4�o���m�@�B�",.�"�G1�ؐ@�\o�����N	���YD�9�1
9���������m�qD��j��eﱗ� �Z� �|X�����B.�/~�}xݵ��q�Q,?�Jq��J�H�p�"�}���q<ta�8���f�ULWJ��U�}\���3r����Ax�C��?�<��A,ou�5�3EVq�Ji�<�R�}�J�8#c��$	uoE\MQ�Jr6\�/9cxnH��0ʮO:I�CT�R��ދ��*,���伒�YI��,вJ���e�x�YP(�|����c�Z^Z%fAz/�TFSy��']9~o��줌�
�M*SE�`8�ۗ6�J6�z�q�Dc :ݼ-��S3X�؂a�a;��8w~�zC@z9S��	�|Iڈ1�����A̎
}����������˹?yӫn��7V6��=��v�h7Z�7���?t�����h�%�Y���Y+����Y�������$�23�l��d`�*彏�,�H�f"p`�`Z9A���֐��&rD{�����Qs�t�8gٖ��f�Ǩ4검��D@*�&|�4Ye0@2В�Bq:�8��"x�D	2��#0�-۽F�(|�l^�@IN*v�Q
�e'	B�Zk8z�:A( &� bE]��nPÐl�?�V�J���HαlF6��y/pAQ�r�g�u��d��x����]�Qm���㑯����,kG׵�4�U]����N1���������T2F�b�ӴY�Z|�#�T��֙3��<�]KO�����np��̺]��V�鰌���Ho�8�O���hѦ0��+�Z�±��Q,U�;��i��p����,�4�T�B;�d\��;2Y�$����!�c�E�]��+�s��	���u�t�9#w�D���A�Z�H8����o����������W�{�(֏>e4D#����"�Uv[0�gGO�kk[8���g����^�B����9x�ŉ��[���)�o���T�K����$�mi&Ֆ�1
9G��T ���]e�eV��5��������%@fa(�;��y�ː��m�J��d���ar^q�D�7�L�)�nT��)X�w����fqB�eY0َK*�,@�5�XC&����Ŋ=;O���}����F��a�s����og����T��qke[C�VI���*�b�a����q\�Bga�7@�>#y;_���:��E� �R&{�E
;Hw���T�B?LT҂�1;�|��p���=�ӹ���?��k���l�o�z_P���Z������!MQ�˂&�8���2�Kڬ�|�Y0͂.f �Ɋv7(3�5u1��mg�ki�����s
���(t8�c3i����\O�G?��G��j�惇ʽ�U��}\Pc*�*&����R�M�6l�OB��V��P�+V�P�v���TC�Ι(�)gH��Lϊt`w4@窺aa8v$`�x0rq�m�9MbI�&sT���vc٩ok�����͇�9�qBe�*(���Y��e9���&LÎ��Tu�_7w�\ES���w����l{I���m�vl�X*
�j�ܩ��êm{�9�OO[N���%d�~�<q�������w�������ƦV����0_-#���lC��$�%Kڿ���/�ַ[�M�A�L����ȡ�((���4J:�	�W�w��ĒToD��2k��(������<w�@K4r�Х�K#{���U�؀��z�@�^C%��c�z3>��7c���8��WQ�M59�d\q�����g�<��owp��C��E��C%oJ���ۇZcF��Kk�����0������b�� ���U�N�
-�)k�+�nv���Bx�IG,A'��o����߹/8?��f!*K�-;�]�b�%Z\DY���OA��	K�eV�,)�Hf�|�,�2���=�ה&�pp����8�:���RV�=1}>��L�I�D���\�8@,6�ӕn�� ����	X��I�����������E8�����>A����;G)�$��:�>qG��Tڕs�"��1�x��� V䢢8���K�ڗ_�?��������v/(�no/�{a�}a�4��h���7�f �����w'�^��gf20�
�W>��Jʑ'�P|.U�>����|��e������ɖ�?�b���<��c�{�gM��>�?���l
}�^Y��ry�
=l�H+��9r�z�0s9�(cH$׃b���TEሁ9�^ɏU$�y�����V�NΠG��!@'�����@��	�l��55��	u$��j�;�c�Q݆z��F�X��(�d�3�<UQȃs�ժ�ku[�B~Ͳ�5�:�en��KӶ�����;y����k�J�O��=���җS�bk���W���{z��iVe�����1R0k\��0���j�z������|�C��8�p�ȕhuzr`�_�'�R����No���,���� f�AG�����N]QjS;}�5��0k��l�]ț�`�N*Q�� jEJog?�������Xy�<�ջq��ð� E-jb�*ZF��ik�p�7Q����L�����}��X|��]������虋���ǡT�;�(��sE"z������g5�c�&m�̨+uH�Y��0�n\�<��Q��Y)�pʤl++bV���t%G�-�&e�_��ZN�q�����sς����r(JA�1V����"�z�&+��<�b���T͊|�R}K|E��6~�h�l%3ւ�+fa)�X5�9U̓9�lЍ����v�v^�`usA,���l"��	����ꧻ�)�����mJ�!$NC�j�3vQׂ��q�������ѭOܦ(��ڷ���v�\�u������������h@�W�Mᡟ�n'��U&!c��N�X'?��@+�A����Nn�ɶ��s�|dc���*��j�V�w�������?~S��ı;�KU���y�}�:���pd��pֲ�;n(�[��`�@#6�)e��"��T�PH��ڂpkŒ���\��i7�#���S<<T��P4��\�<�3Q���:�#��$s���-Dj�RT�|��^��
�5M�5u���5���i�׫��J���v�Z�,..�u]w��m4A�P��	Jz)���坅����ړ�Ӈ��"Nnqn�������� 9S�T���47N�S���8��/��(�:��ƾE�v����ګ�`"�U������]:է��1�j�(5dV�%mc�l���.�7�!��I����C�Ab
�wyg?������
���/p���p�+a���@��M%��<u�;N4����������6X"b7�Z�����y�{|A~cй'U���D26r��e�Ny[�a���^���q&�3�j�)��Y¥�����>A
d��o�jHj��f�h]ը�,�)zIM�T��Oe�90�.�C�3{O�~B��2lJ����)�"��	Zy���AQ�!�8V�i �*�t&D�
ι�%4:�ᰲf����!o�(X:�<�MWQ+��ä���`氺�%�Y���f+�FD�����1	g��ua.d�A|s��*���_{�GI�?p�b������=7��A�[�����2I�����ﻴ���V2�M�}rٌ#[0��\�{�-�����-��:���f�u�'j��&U���'�"qq�bL
��cF8[���������]w���WjG�ַ�k���m���j6�7�7�o�l/���"0�ʄ���R[áT��(���z.
33�N�|�B1����Xi�
y��2��%��^(��l܄s���6��0����D�c%#j8&�]�qM;7Ve�hZж"��5˶�y��i�;������Qa�<V-˫�7���k�.w���_��?~���Ov����n��KM=����W����#�����@��?���p~��ӫ-<��q�n�Q�M�d��✈7�O2?Q�����`�A��ߗi/��T~t��Z�՘�΂`Nm�!'�͋b��vB��^VX4}V#��uԃ.~�G?�w�v-���g�]:�z�=�Q��T�u,{���*�v\�n�E�jfjX������cim�Q �~ ]cG7|���������Ô�j؈TZEDY���N=팗:�=K;�Ed��/;7�Ҁ%z�v*�Έݟ|,XS��ܑx��j�djI�>J����	�1�K7�|}AB�1��2�r,0��#H��W���19���xlYa�r���,Kj�	s�-)u*f �?r��x�1��wM�U�߁ҫ�GA�`�!n��*����`���^[�&die����kh�cʠx�!��>E0�vr�Ts�\`9K��>x    IDAT�T��>j��#ӥG��_�\���mw4^�����~�F��Zz���,�����q� pg�-�N��w�:��v�l���ߋ����LJ8�#�KU��lw2X�aA_rf�&�%n`K��œ��9jq�w�Z.|j��[�rM��Gsu=���6��a{��z�ѣG?��tl�
MF�
��\�j5�n�HH������w�Պ�;�ڋ��l`.Xn:q�B|����#�+��<|��%�P��8*��nR�F�XUAt�(���p��ϟ�usm�:�<=;��(��Rn455�������C�R���t��V����k�8���Jn��f}�2�T<y�,�>s�VO�g���h~������~�}�i,o�pag��=�,B7���Z.	h)��@I�� [�.,��e�8H]�����"��T�H-~��sD@>-�O�d�9�?U��3oH��tQ*Z*�K��Ou�+?����+�ȟ��=ʖ���x���m��>�|�-��Lk �h�ĵ��0]�����|��p�x�F�+�<�amh�(5�EK�]D�#H�ؠ�$���=E�+�-�p���L�%8�I������2R1�J�`��3�1��3��"#��ن���XY�.�6L�5&F���U�K���8e���U�w7p�]��h��{� ~�9I���{/�X��$����D����]3��Yu�J �$f�G�s��"T:n��F�J�4bn����>�~rK#;#V�#i'�L�#U�5i����]��.�D3��RCU:<e���W6���\����PA|o�����#��&[������&mV�
%�|NY`̼p�G�͙�ei�F$9S�	�i������{F+:N�t��'g�H�H�G2B�}��Q8c����R^(߃�]C���_W��t�57?���;g#���^��p����'�>�kkw���Y	�}"	i�V��LC�������(�M�@�m��I4W`ц�f��OZ�!�	�
B��Hӵ�`����7�]GU��x�l���E�j�VY�V*���j�T�O�-�f��b�QX��H��F�K���Go[m�S�/��Ss�R��'�p��9l촓9&u����M|��o��u'�����c'������O�3�E<����L�
MX��2�� v�]�9iA%��k(S�n���z�"Q��5�`,�H�Q�m�߆��0��k$�:�Y���c�zG*�����vx���_j����t�7�� .�p�=�_mt�T{��͡(�Wr���j9V���б��@S���r6�
��0K��#��ܤs��W��[>�fJ�#�'��pd2K��zA�8I��H�F��R���"��i����]m�(��R/�NQ�yǋ�UH"�Ϛ�5�J�}���K�O#�9+ʉDYȌ֘���&���ńB��r@^l����3f&�d�!@I�:�&��V���Z����q2��#�N����T����`��ը`�i��f�6��`\�<h�S6	�Bs�U	��0d��h��,?�\�n/?r�5�~�w�u��|K�9^PE�E��tj���^���a迂^����,{�2�Ƀp2pHF<�j6�@��]p�&n���g��"�K�\��e!Z3�ͼ}�S�D2ʀ$���'4
(��p��� ��8�{�㸝��}��	���Ǯ�W�l��(�vЯ��}��(
Hg7�@bp@u�^�����}g�%̿5J~�B�����D"��3��#��s��(q<��h��F��nl�J��\�d�Z�(�ʃ�����}���)������K!(}+���3�W[o8�����P����Wڎ���]���(KԼ°��F����y�C����SKX�v��=�����jA�&�S�ZE����s-p�D���J%�$؄�P2#�A4z�Vo���$��CЍ<W,I�1�&�F����1���m������3�}	�;ā�����f�8e����>����8~~C(hs�*�ZX�s�P��1v�����3�졗�L�¦[F_��(6Q�W��V�O(�*ŀ��Jjls�E��n��ِx��$���,=�}�V��"�|<Kv�&�IU��(��$XK��e�5�{�$�i��S�1?|J0f4A��bD�t�h�z��疤b��� M�ҙ�@2�Ks�fa���Ů��`�!�6�����=2��n�K�|?I�=�����k�p������5���>y��UXn:����ن�e f�~b2��Q̳�N��@��R����`��=y�l��,�_�i߾oɳ��8^�u:��a�'��{s��dF�Q��;93�*[��鎜�[2�s�h% 1;���Nޗ�����JYn�&~�B��M����t�3��m813��b�����}�?�{���_�^�mo� ��f���pj0v�
G�r%��s`PBDA"��\�{�szv^@$�]V$�<ʬ\�~�E�u�󼑦�tl��k*Z�N{�X(��W�'����l��(����T��C����坊�;�����N���q��G��x�kOa����wy}���y�����ڸ��'�䦰݋pa��s��(��*Қ�l#)��þ8�t;=LM/���%\p�	Rp%�E8c�'d3�����H"դ9��Jf�)z��X������2��������~���<�0�1=��mà/*�ߊ�W��%��:��^��GX�5p��*59��>6�]^���k�ΠOa�Mc��r��'�Z*F%|�DQ�5h"8��x`�:.���x7�^"x��*q\�όI5��I�Fd3�,���l�3в5����	�S�.'��D��߳q;Y�\����&���r�6yNv�&���l��zRА�ȱ�$�1[��!:�\6)�>�����#�1t�=�Y,����cy��J�X�j�ЧL,���AU�f�r�r!'�S���|���kڧ_~(��3��P�8����l��8��}��QU^H�eŚ��0�N�a����^��Mɺ�mc�=+�T<"����a��l�X�J�(�x>��?�������:��~��wr�b=
��̾iskk�A*��$�saq���*�#����%:�[L����'�Ss=���a8�A�QU���z3��%�4�][�T+
y�����^�Q����.����륞qygg��N��g�ݏ�X_׋�8�����u�,/K��������x;z��}�)�Z;���oce�#�y�z�@�@����/I�p0�����$Z�iۑv�\��bC2���"7�3�0tU��`N�*�Q4
���W��܌��'߃����݂�$*cEÀ>�1A��mn�;[X���g��X�s�bnuӆ�X��;P"��~����YCa!����$ &z�|,�Y�� �(���p�'΋L1���c�f�?&�!�g��^�e��l6O�7.%�N��ʙ	4�U2�Jzf�P3��I��I��('��$Ͼ����&��ū0ІToRb�J-�+PA����f��@���_Tq�5p��y�9l����l����E�	1��s/����0 E�3Q�
F(�,��@��Z�=Gj�nڟ�r���7��n]9���G�0�'f�i���e����!�&�m'��'����-�L�"��\���2�� {���=>�O�wI�)��8y�L��O�˥Q��,{���6хGTW�DT�'��j�\Ŝ��& ������9LZQoT����+j�V)W�J��3�3�K��v}j�?]�]s����x�7���K#��[�Vqs=~ͅ���_?�|��H5N]�A`��������:|�ߎ��-|�'�������Z�:taR�"��b��O�h�Q�vR3���9�Ĥ-[�Y%��AŶ�O���#�����64���r�� BpTN`�=X�5�������[��_~�aѰ#�q��u)R���Exlg�c{'�c�[�#����}��=��uw��=���
��a�Y�iDv	��"�%hy�9��ka��-��3$/�LŕjR�5�;d{������H����=ۿ�� ��Y)o+���5#~�q�����ɕ��GV�&#�g
Vd ��~{����r�b�")��vY'�يy��W��`� 33]&!� ~�t뒛���������x��W���� �N�z8����V����Ǌ8��S�Z(+J���� �9mшp�t%�1�{��D�zف�×�%Χ�p{�q���8���~pEF����6��-��lQLҁ�2B��/�)
�-�g�{�ϓ��U�,~�u	 ɀ)�Nt��e��&��_�T���ja�⢽��������u%��$���������D�.�.f��mc�����Dg,>4]�}>_,����h�7M�X�~K���燾��g�RԹ���V�ч�X꼿��˛=�F>�?}kK��x�;��z�p��I���Q<qj��&�7�"�D�Ӆ�VB�\��Ѥ9;Q�Pe�@��1O�|������H��i����2e �]�zŲд��Z��i���� �"?�į���UU���(�ȅ.ry� Gl�fa}�������'w:������Ç�8�@�E�t�a�j8|�:��z��aݸ��,���Lq�y蚍 z"X!�61`%�@�����K�,��QT��u/�|$3 �)h2"G��G�B�X�8�N��L�/>FP�͑o��jN��T�l��s�� ���j�X�"N���8��M~�g�(�	�:��j��6�6�%Ъb��!�� �E��^}d-8���gW��w1��a@G0���KX:{�a���=sJz�+��є��s��O������%�*��p�&����73Pf�������hS��tN;��@;�j��p��=�:%(�	��ɗ�;��,�\3��%��3�D2���B�#�*5������w��n�;-x�	�� �1n(�{y�Q����N���r�3oVD:�02c�����k�������[���d@{��M�	��ܜ���[�?z�'�v���p~iO=u�N�B�R���>��U����'�ı���'��YF�ԐN
�T�ZA�R�댰��-�jqTI�>�<���
�a��Q�VT�G��L؏�Y>( AT/+9Ҁ(f�����8b���?�C�t�|�k��#4r���|'��]E��>�l��p���:CO `7>��j^��֠�V���LT��1��h��G#��@�u�/�?�%3�N&�:ylCRk�e�*����Z�Ypnm�X����Υ�aZ�J�� ��M��?*�)v^����.�$0Dr_L��`��c)Ň��re*�:�/���w3d�6�h�$~r�{��3�'Z���!�x��T�J�0u�G�Hf�=��v�0���<��]w%�w:8�����1���)&�H�Q(c�r��J�{Φ�����@��F!�6�{�O_��r�mlll;|u�����~��ifV��#̄ĳei�>�q��dv6Y�^*��jLFH�t�I�I�\br�f��-HɄSK-1dNeڈRf�K��\_��>|�g>��}s��TС�cG4��b ��J� '(�(:�t\l�s����3�}S��������=�����o��r��~�v�������'�8��Qh࡯=���-��.���}�H;����Q�m�{�fσnW��e��S1�C����K�'�#�Ů��1U6�V0[Ɖ��qƉ��|.[��U^2㣴^DN:�5� �!w����Q���+��w�S_G��Q�m�,9[G�ۇj��������8�xjs#�]JE\{`���Q���3D�f�t�R*�K��s�U��"�>`z6k������&*@�{�� ��H���&���mh��P
0�J�N��e�qʊv��Jxw��\��>��T��$kI:ZI�e�4�$�y���U��zg�6�3�}�2;� ~Q�j�����DE�}��Iǥ����a��0����I��W��œ��M�Vt�a�w�A��뱼����6�,�a,��yx����@/���Qbh�)�R������V�����h��F��v�rE{�#4����^�����C��~����@���&I�@���Z��&� ���2��q.��贓d�{��h��sLV����I��!sE j�)����Q����hm7�����kw�G
|U��l1��?�Z*�������!��I'�u��hҚ�*���
U��8���L7���n���K�<y9f}sq['�wn��Ǘv:߳����_�ò�lᕷ���5 ������ ���'��u��H5�:��K�~�A���<inb�m%�, 0Hp�y��#�SCAʦ8
����E�_�n�
R/?R�G��(�m�υx����m7_����l�G-1W)�P�N�	P
�,��V'zo���sh��I��r~ESE��F���p�~��kXs�U�:b2��s�K�ea��c�؅�klN
0f��${��������$��Q/+��K@k<�F*�1+k�k���T<i�P	6K���,�k�4H��������k}2�^S=�F�y�sD:pi2��u���wϹ�2�W���@�\I�jy>QPG��휬3V���	���x��-�^�o��*�<���N�7$�JE�q ��$�-(�.�UT
t�w�!�x��Q���#��_�p�~�r���gQ���u���=����A0ÛM�V3��$O$��g�?s�y��*�/u��=�3���.���MJ�K���������������8wꌈ�VAھ�k˘��0춥R-�*X��D�1����e{��Oc?q�I7���9��Zܿ�KoxÝ��u���'�q�m�AN/tA�����^��?�kx��cՓ��
R�k��oz#����gVv��׏���K�:J�}(�����c{sC��t�au�o�2��Y�Z�������9������	� �p���2K5�Ţ�]�q�7B�N[�oY����~*�Ml|�̛�6�P/��Q��ac'Rp��n���������,�a�Ra&�4�pHqӊ�5� ��a�T�vM��T+9�I���0���}�d�r�J!v�(!y	�Rv���gd�#��1�����V>/�c�ϯ�T�*tE�<�`�ƽ/��Ԏ�gC꽓>u�	!�8+���%ۀ~��#���Ln2HN�ä���a��4�pdT������3��R��ͺ*�x�ě;g�EK<~��^~���Hć��k�>�Rm
�W6q��:��YD��f�w1�D��O�8�i�WkKE{E�M[�{�(�ӗ�s^���a���5>�������)���l�v�5r���jn�v�~�@�l/}��If�[3��xZ)��:i`J9W�������W�a�^��,���\�.�'��g�'�1bk0Ā��R�r�AM��v��Y����_}�o��ͯ��G�k�%+.���	4��ť���T��Q�X=�������}3��?�GNl��fG�,ai�O�#_��mj[wZ;������A�[�F9F�������{z����A-���*[�H�aǆ#B���ߢř!�jC�P6"��m�;��;oƇ��P��b��G��hCQ4�3�;;6]���'/`-�ql����CՑ��Q˙�����Fez�^�Ȭ�h��������&���������fU��x��>�锝�~�E�ĽI��rS���׸ۂ��]'�p����lfYK��V4�3��+�?���-O� Mc�`����j�G&`(��S�����	�����b��u��.^���v��� �ŒoRf���ޱY��{�c���m�"�D����]�5~sSP�?��o��N��ⱧN@���h1
b�BF�$�>�褓B�h�?2+d;�p�t)&��H)����.W��r����3|�x�~���k��59;جu�eW٢yg��g<_E�w6�w�=��i��ٮ8��ʒ��c�B;�x���U��[G�
��r>'�PV�W\��V�>�V����N�]�6��1/�rim����_��;~��o{�S��v�ed�Y/��nl�g֚;߻�l��u7�z]4���Z**�g��Wp~���˛��ᱢ3���D��ԛ^��^�%�����     IDATm�Q�T�*:���8h��fV���:=B�*�l͓�J���QP�!��լ���8��1ʪs�}�>����^����\8��REU�x�O����-�e&{l���3�h��V�ko�N,ڊ��lv{0�u�<Յ�����9���Ql�ﰍ�XwR��B۰se�,[A�$�^B��j�~�-��Lv﬒����a
�i2���J��25�y=+�T�����O�H&��e��Τ��$V��=lL��/g-��6)c�� -a5(�sYj�29ۻ&Ͽ�A9�$Iw��C���.B�r���V��*GE.J�)�)�����q���/v����k;�f#W���|֤)AW�(B1o�F��p�t����o>�{�2��Y�f�Y���w���Ӟ����A˥/�%`�l!��'��/�l�f�cq�-�竈�$���S��0�(/y�!l�D������g�����z�XF莱�~T��h8���ß�� �^�!�Xۖ���4�6t����x�Ϳ������|�{�se�b�K���;�7>~��/�[<p�)K�va!_Bl���u�������]^d�Wt8n�ʅ�TN�NK�a�zcF�"��&�*�v��".Nn"l�ʖ����J�Lٚ6,���O)�(�E9 7\���:>�7�1ncp�8�~W�l)����&J�2�q��(���.�j��zK���㆛nH(:����5�Y��*��
<�Ǯ#?{vu�����d 	T�r]~��.L���ϠbT��mJ�g\4�\|�Y��l�6f���
�<WRo2&B�.N۽�C�ȹe��b�%0+��S� %����'��d���5+iv���#�&U����$�"��tH
����	�d`�0J��)N��.8�g���̖J���苼l��	h�T� S�"n��F�P���-�f�J#7�1r�M����#�Q�Ŋ<�{0c��.ş��`��ˁ�Y�8>e���m��}�u���<�4�5�4Cy�u�(�dA�u�T5���g=�=2)��\��t�)mf�E�X�ż	�3)<F�V*� )@ֿ���s����4d-�|�������Rr�Wp��Sh�Gk(�N�Vq$�pζV��o�����c/�8q���O >�+v�U�Ϟ��k��k�r&
��\ĉ�8��ƅ�.V7��C�1Q�D�&X�`+���GX]Y�6o�\������k�h@g{Yr����kkk����Rڛ�Y�b�]��+�9(*c����~�;n��܇񙧠t6QU5���K�i��w��BO��xd������ 6a�󘞟�\�����`M�#4*����rthS��Wf��g0�� �M�rǈ(7�w�j9�|�UF�ׅ�S�=�,��2���_6_}�s#q�I�M����ce]8�����j�6-����/bF@�-jH+�g&�\��� gӲ$�3�&4�d6�]x�V��\�?3�xV��3�ȕ��4	zY��7�f����.D��=-�\4 ���'
��
����l�爡����~�k�ؓ�X����v��9l��ȗ���:���=�3ڜ��c��cE�իJѧ�(��������v/ɻ�`���w��s��8�{<���x��˲1.�D�b�?���/�s�-YxZǗz�l�Q�-Y�i�O	�98�%h!%Ж,�����6~����*�)8�ș<���"6�>��/�<�����$вm��Z�M�h�O����~�u�{�_\�f_�:x)�;�c��J������SKko����5�΋ŗ�y�#[��[C��H�#M�{�wț��j�w}mS��֧�>�h�NY&��n��Z���I�ɀ�� �,�b�a����Ù���dƨ����E��O��m���?�R8FY3��t��K��B�(��V'�ܳ����Jl`~a�Sp;+K�U������毿�U����/�:�BO-�B�W��U�0q�u��"�h=�hB�8���]e�c2/���mt5Q��ڨ��?����51[�?�0H>g%B���ؔ<�"�V�A����:6�9��Cf~�ҢM=c3C����e�6�^�R��1m"8��h���nҐ5��|��^�1	 ş�T���4s%���;�#J= O�?���ѣO�]�������pvy�r��+Y�Ը�h�`q��l���v��+*ʿ�f���mWԻ/Ž�b_��I��ύ��.��~�u��|�W2�}�I��M�v�Q��h�ǾT�ǿ�>y����}���*�&���H9�x�����?�R����������<f���X<��V���|me�@T(@�'m�Ա8U[��M}��;_�[��ǎ*ʄ�Ջ�@.����	з���k79q�s�P}Kh�JF��Vo���m}�4"3���3�Ev�;��x��	�@)���Q�ǥ�,tv� -�XD��&ʘ5��i\�m��������t\�v����������C���n�G�|�ӏAo��80"��@���T}z.�;8����
����l�V�ajj
��"o����
\��Ȟ�n̢�[���8jA���w*Q��޻��ZHM8�	Eˡ?BW�h#*�6BzԦ�݀�V��)��cB>��
�#5!݅�f�X,�b���Kj��9�:P����i���W��n����|r�$�$�7n�ٮ�x���Y����dk8K�����,�NV���0y�f�e�mLg�������e��̈́�ϝ�mI�l])٩Z�n+k�Jk��]���E4;}����!l���iH]hq:
`�*����a�da֎￪�|��F��ˁ�9N�V�L%��;|�����y�����6qV��!2_����~1
V_���R�	.L���%��|ErZq�jŲT�4���6�V����_�O|�sx�u�asi	�F�RG��a�s�$~�3��jñ��JE�y��\yh�����{��]�y�[޲�b>���}�~[����~V�*���u��׶�8v�r�6�=	0#WA�7$�R���R�Dz�.z݁لW��+�x�Z4���M�X<f1ug���݇�sS[=�}B�g�����0�ҏ6�@���+��w܆[J1���(AY��T]��ȏ��*v<����;�����Q� W�-ʱ�r��h�y
��"���b�0��<��<FZN�3�2�Р�<�F�&m������D#�P�ܮS�$u0qy���0a���l�*NZJ,�B�g�BqI�ӥ��P[�6�ݎf�@��Ң�hw(�*�s9�A(�+��L�-`zn^:<�X͆�3&�7m��'e"\b	gc�Dn9�`��Di��K%�Z񩩁��S�]+I ��<$O�	ix.�DF�l��P��f+\Zٮ+�S��t�<����\z���M�x��p�����[q�$����ժ�G҄꣱�����-V8�b5�9;���i㗯���h��,��sv�k�,�÷���:�3�@ʃb�';�IgYU�^�Q�ҿ����X��6�$�fIKU�D�=L���A,H�����#2eE��W*�Zm|�O�'��Q�b�M�a�9��7�W���ş�� �b~��Z�"�p j^�u�W��{��o{�2���~�/���������|���U�[�����`u��XC���X�n�u!V�T#j�A�@<V�����n�����,����Ŕu( ���=.�2LUE��Do0Y=po�D0>� ���\4��_�[���O����>y��S��!4��f��\En���~�m�h�7{xr����j�Fq���D(�"�C�R�]?�О�>}Ae?F���^�=2�}��Ll��s5�p�_�xFҢ�T
�����g�A���jI(Rk΢^���+K������R1%�����n��\����<�j���.���9��Q.�Z[�����r���YUM>c:��|�+E˥,,MD��%�|)���{6���+OR�h��5@j����>�F��)�����w��a������x{
p$�N2��JyW�9I�:y�M��&iK-v�X��L�x˛^����+n��V\X����Alt�H��gh�JW�"��WQ��֜{o?X�������i���َ�8��nw�H�w���u�*~A�{�3m����=����C��O���٢�|��:E��%���2cf6-vW
��)��X�be�:��Ӂ��V����RbqfV�Q���k�ï���g|A����#o٨U�0����O�t�-��u��������g��..���	lo�Fݻ<=���Zm���e��{��u�
ڽ1��1�#c�����lң��7*��h��AU��z�!LB�4N��PL��\>q�	��6�L��C^�fR�[;=��dP�>��&n���]��ǝ�E4��� ű�?t�G�>�A�,����C<����Ϭb3TQ^�G�Z������<<��q�YGT]Ĩ0#ڸ܋���)��xr}��m�z��k���5�e@��.Z[�tvĮ-Q�
E���t�6�����^-�aU���JJ.� ��!
j�\8Fk��76Иߏ��l".����5W_w��Y�H��8SO:g��Fh%�r����p	F�-[�N�HXe��lI�IyH{�l�fD��
a[���3��L+>�n{ =�,%��b�{�(,�,3�"�^W]u�/�cih9�A�q�n�.�Y[Q�l�)�ǌ2����_����{�/��>j���iߏ�p��'g�jEQ��öT'-�R@e���	��wN�l1e�W7r�SG �\Q�a;Zf�����ֹ�gƳպ7_i�[��PG#L
x�/�;V�:���DQ�z�mv~���O�icd0�	�Q��ѻS������W��;n���7����{������	�ٵ��C�?�i�+�>έ툫��+cm�����vp�7Ā�f�4��d�v�5�@kZE9�x��x��e����$#��Ǩ�A��#���@t��XVrS9�%4@�h��"?��{��V�����'�9�+�6���%4��Á������n���x��>��������PM���\�6�m��jku���5xv�͋6./�'S�V���U)p2qf<�1���$��i !��1��x�H���Ơ�-<ND���K�2����(�R�I7`n�1���:��	��D���Gs���WP����¼Ш��{���ȕʨ��C�RÐ����%3�& �I�����d�+s�=��}R��MO��ǝ��x���$l���*�.���:�}(���<�|�b���]/��x�C�a��Z#�>}=7�&��9CE��T�s���+�W���6J�w�?�+�;C����������G�y'�r&[���0����*���O�u�7�v���� �C7�C1�r��=UU�M���a<U(\���5�-�&/v{��Ϣ�����0�1tT`��ԇ��ʯ����!U�L<E)_/�V<��;^�o������|[���M�	��������F��qW����6:Cl4{�a�鳫p1��c��#Q�aKT �i%�F*���vzh)���s,A�3B�0P����\�q ��T�!��@�@C��	WRCA�����`/���7݆�U����A��b!g!����H�.bE!�Z��`��������v�
������7�����3+����1�  H�(Q�HQ�u��V[��v�[�J\���5%�nY�h��k������k�hZ/�	� H` 0�tO��uW�}m��U3=C$@�8:#:z���*3++����,�j�Z����l��؜��T�)Ef�!$��+F��r6hw۵N��&M`����ɡ�3�gZ��P�L�-l�.CS��{�Z�Թ�9(#>*���ϣ0Ama��ŋ�$���R���XAw{�F��<b�
<y��G��\A,�D���'tcY)���Ԧ��?�Ԧ;�*��,�2��:�V�[Ez�)_��v���V�S���S�ݽ��5-��vpp�������� �>�3J�?���%�Y�R�&��D�3���|�΅���V���^E�76bXvƛG#7�1��~>I�����WV��?�u���*�^a=�n�Z�Ǒ@ϋ��N�!�����*�
~$H²$*�i���?~<�i�Q3��q��/�ҩ��X�qΦ3� F���a��ٟ`+05���@�7�d�Q{���7��o~�'�HP��|	�9k����v"��'h�Py�y���M+�e�*�k3�l�b�zl�������v;}lm��������ļ̀9cؒv�4�"K)��Dm?���^ ;�P�#h���`+���{	3�|�Mx��9(��+gАE$�r�k:�Ut\;x�qprc'/-#1�?z�����6����	{�A�
�"�B	��@h� ֋0is�lp���L7vWX��[���@���r�V��x�����d!8����bY	�p��9>I:?��ǙƝf�"�T��P�yh��m��w�� �$@k���(���ڦ�����(TjRV��H��
/nxr:�f�uL-d�j ��2�}O#���z��J(�� �^�\����ٻ����5���f݂$[��N6n;'��Eظ���tx	i�cqQ���O�������1��0o���2�<m^Ì������T��h��߷������fDϿ������qQ����s����纗���n���1�p�0A�>�d�O:��(
۩ mǉ���B[�#7�}/MW��b�/	i��j�ɬ?�W�T!m_8'|�s�E�H�*�������#I��?�tT���R,!��0m�87����|�{��zω�K���=�Up��auk��I��x�|;�IG^���-lw�x��e�Ղ|��2t����֕�� ��.67w��8g�����Zt����	��H[K��a@Qz� I�S(7�1if�%N��A�_ĝ�:��=�`	.F�D��q���&ˀ��0���܈xt�2�
2�|�ֺ=�Q���б�z#v�"�p�M %xb#���XFb�B-6���t��w7�ҿww��^�v��Y� �D�\�+�^�$���3��c8�YD!�s";�2FN�.[H�҉�!Ɍ(Āf������8�	�4��� �G@� B�J��n����f��W�jM&SM���6i�L�U�6�reM|���]W�ܢ��$�Mg�\�^�[��k�s�+ħ�L6=�S9�n�*�n���g�dX1�霜*Z��\0P+��,�p��I�����N7�#'Oa
�� k�(�GQ0d�ݛ+�˥��s_�������7qS�|ZY��A`��a�� �5����m��������yf�tuF�(z D#J��~�	\@&I∢�!IhA�j��/��v�� �
<��9���������)����o���ڬ�o�׷>��q��fv/\���9���b!�@�D��`���+�/`�h[�è�Xir�����x��o��}�{NP��5�j�����:��9�������@mɍ�6��<yb�͠�VCo�b��lX1%�d�t�ln�e,ô��쒨��BġI��I�[z�S[�n�@�?���^�($@MC�>n*x��Y�3�Aڸ�x}uCǰ?���ˁ�c�� �3�pql㾝.�jqx �(��;#6x`�� A�(P����\Ŏ�s�8_������U3���,���'��'��9�l4A��R���	���h��-@(m�ݜ2��f��x�(
P.W�RyO1{�@v~-�%�(	�T9]�
N%W$"�>9������:��j�n�<���4&���g,e��	���*�l{�K`ZYN�On�RU+gd����$������2 �� �V�q^���=+�^S�+	FFx��=EK�?�Ab:m��~
����v�[]�)�;ʀ��M��Ʀ�jN¬�`��}�R���C{@�M��(6���\�<�(�?��$IE �n�������^�tiG��r�I=�y<i6/����
��t�$��T�[m k�<$R�$�Nʾ����iA���J��&����k�������`������DpR��3���ntDv(���aH-    IDAT�����/�DVř&������c�n����y۟���{6������W�X��ˉ��ү�m�n���D�5���A"�P����t�t�'�����"!��n��@+�*
�
G9:d�O� q6�%Z/"�P:�O���ΖHW�md�,���6��:~�>���h/�9s:e�
�X�Y�����1���1.���� 㓫�X�<&U�l�[��-���Fz�D)@-�c0�X$���Y6�'�mS���:u�����p-j���B��P&���DA���gg�E @�N�<����I�,Ѹ�# ^,��4��L�N�B���#q8{�i�8q��]��c�a�!$����m�:�ç��i]���i߿dwW��j4`�C���9�8,��S}.�NL�;�CӪujt���A����W�6$�C԰�B9��L��c����U����/�S����ːPʛhX
jj�/ȟz�B�,Y7����7u�[]]5r9� ��9���MH)�<\����W<hHA���E��-�(IҎ ��4%6�	)U�^���$��4��$�vKAɁ��Q�&I���P	�C!˶zQ-�'��{����\���K���8�aaf��0�)
�.{��2~��#��TCyv�?�E�<�����>�7?����^���=�Uu��n������^"�)L$ɍ ۏ���_}��e���\o�5�&p��n�;�z��60�!�:	Y9F�W7u��!R߆A��(�%f*��fYl"0��2�
D豋�����'�|'
1�3���h��GR0)?V�f�?¥K+8���w���`�P�\�R�T�Ta�F�P�#�a+U��\D��D��g�) L5���(�*�+��ٹN��ڤ��̙IU����mb�H�JsZ
� ��*����B��Jwnn�^"'�����8|�z����gڳm��R%L&�b�����@Jɨ�C�QG�3���(H���H�5�NH�#�l�H�`2� ��\��W۳�U��I���������n���jz*9��/phN��)�k�G-d�����&c������{S`YPҹSɶ�P���=oj�>y�L�_2�G*aς��������k
�$-i!�e8K��J�4M�6G�S�����K�0M�~F_�*�X��8
u]��$��4N�(A5�M�����r�S�*�~����:���۾QQ�[�כ�^$��11-ED�*>�'�
q���ðu�M+)�/�����[33����PE�����@��+������ ��B��0a��q,�� ��av� �H����c/�3��x"?��j�'��I��d���=@�;08��ؠ?>��e���u;�0�1������gA�<c�,�3J�]�AD	|��s}lu��p~�}��S���u�3�j�Z��w�3�b֑��(��
�:��W2�/�Q-[�_'�̜��9�T3Kև�g�Tk��h���bH�f�V2� ob��$9Q˘Zġ�a��E���9��ks������mK��߾,q&�6��+cjc3�
)�B	�x��s�8�a�P)/XR`r��j������3kC2� �,�2r�����aZIO�yw�����kj�O+����Yt:���vm�����ny�R���r������_{;�>ƮQ18��M�D'-s�`�aI���z������r����k��m%C�>Ai�*�n�PW�l�"����z*�@����i)kR�-��،�(�����d����ײ��D��j�=�Л.>�����w��OZx�^�Q��=���~�_�9N����pb.�F��K��������Fy/w���~7^�������D|S"H"�H/��O��(P�Ρo��l��G��HP�*��v�����"���)Y&�!��H�e=\�Q?�\�d��K�4�7��نب�>��h��f0���㘅˳����(CΕЍt��b��q~}g/�`��`*0�5(9W���%�o7pi}fe�R�8�Ñ��2���@Р�&j���h�}���(ɩ���R�f�Ϋ%�N�\qLʀ6�)��l��!�7�a�4T�E��=ny)gg��m4juJ��@M*�4�,1�u�����L��4�:Y��>j�
�-ZV�� ��y�g��!&R�$���	W���<G2%�']կN�
�=�d�������,l��ݥ��4#���+�(Z�L�'��Ud�=�Yˀ�؈7[hA�N��D����Nf@��CĲJ1����Y��ni�>}b&���9����~7nS��פ��}��7��̽��;�5Y2)\��lN��<js勐fg������m��t�(D�Y�����{��x�3��#�ۓ��PE�=��5t�_�T�� ��6��8��G�	�%l��l`A$��Of �7.�&� kT��Ȱ�4����\u�TY�Y��V֑���(§����C����&��#e?x�>Ԣ>�a��GSJ ��� �b�T�����^��Ro���=��V����B������3�yj����0���%�R�T@��

�Tf`����l55T���Y'ˮr׆ \��t+�`��M����D�DjiZ&�+F:X>��PT�Y��![뗰�����"�J����|����n������KP��U�:�R�Ȉ$Dd�O�)E����e���zZ
 �����ȕ�O�_��u8�\��j��W�`֤���g����L�N�%�H��k�&!�����x@�/����I@�6�v�Q��m�w�76u(d���GݿJ��ق��!���m���2܇�����J�;=y���������G>�`y)��/�Xc�S%�Ԗ�s@��?��}x��2�u76�=4��'n�������쮻��*9��|�g�B�[������hSQ�hv��T�z���Ї�Z�h���MF�W���%��x��,4��L
kO�j2�,�����銎�"�D@UD��ׅ�[E5�q�lw,���":g�����QF��df^�T��q
G�q����;x��xD��Q���У`�z���>x�H�
Z��X�#P�D��c?f��ѝ�4�T11�H���,#�t��Y��5�ӷE�TfU�^Z��Y��j��I��K�ry��<��YDl���O��o?�BJ.Ϥ���
����G�:�t�r�"�A,�%5#�s8%�n�� ���9�Q�<�m9o2הhbF@K�T!cx&�,��@{岛�~C�;�,���	�<���)$b�6mO��b�2E7^��SYb�QmTYFy쎵oi�;*�;m��1����)ۛ�ʺ,�Z)���1����F�3'f���/�f�Zyxz�|����/<y�}?;g��jB�Y���C!��f,�@��������s��]X�i�^-��������?���˯�s�w����v������D�;9L(K5��HX�h|HZ�.ov��C�4�iS��\^YC���h%j[�Ej���gȕ�HQsb��mI�L�@���l�hA���q�i�8ڄ��M6��
z�.�u�F�]�փ�(c	��_���6pj��YG~v���#S�D�9� py��Q�B).���*"�_йZ'/`��k�V-²țY�y*U�4���mqwIg�m���(�5I)6q� MQn�˒!a?�|NExX�t�,.d,䂡b�������\: %_�F)YƓ�}傉�f�0Ν�Q(`��qn�S������#I�@�l69��X�b�;`�/���B�ݚ).�B≼�F�Ё]���P�� в���l��Ta�����r�dS�%�-J�!������Z�m&66����,�9,��9n�Z������eh*��f@[�	����M��go���u�{d��;*�ι������o�C��F��(F�R�I�	��y�����SO�Z<��pD3�����ә��_��-o�x�\O�Vj���;�c�#~��-�$���ڎ~*����;���:#�_�a��:��REK7�)�v�=���D9˄�4A���lҘƁ2D̀�aÖw�d����C���fM�R7�O��l��Q���DT����
��E��	���n�3�ז�pr����Al4�Wʜ(d�&
�U��A� &KxI�Lm�<|R��
�,@���z��R�� I~�S$��S�45�a`��obDq��D����Z��`V�,;���cߗ��k�`�
�f��=�/�9�֖3�C��P��A_�x�5�G�y�{���Pr��݊a��A��Q�Ru��EN[���<�b�TJ0�,8�|�B�Y(zdc��u<����������)�O� �D3�	�+�	z:3���Oh��5y}٦a��U��[�IKK�����0�]��m~�r���Ӥ���K(�f�$��i~����'�s�{^ǯ���fz�歯����?����A��\fH�G@��!Fq����x|��{O>� _F?�`����e��}�����;���3p)M�d�wgw0�'~��#���q�,Y���c�KFdy��G8����G���%�&H�g�buu���cv���4��ĮˌV��H
�����t|�io��x�b���6��� �掃\����<W���5
&z�~���/�t���C��l�@H��a���Y�w{#�^ɪ�K�vd�}�4�59sVTT�����x�r!�j�̏'����u-3���+U�Ur�mp� �d��8A@at�'��������c��;(�+�6��/F	lǃU����d��0�!�)��6����3�p���o��H@.��}&e�,y����"_,suOl[z�	�h�(lG��jI����$���乞yA�x ���G<��Y'�rbp!d-݉��՟f����䕽�����>���!����|,3��e�N\�)�Ж�p��GC�P��7�;�s��T�d�0��1�(G�/I�je�`̥эM�3'�����B^���?J��=�������{����Z(ձ;��?Y�Y�"��1��y�U���BP��k.a���������h������*���唦���ݽc���X�����6&�O�]���4��b��ak�p�GLc]��v�����P�Pn.�<P�����ihpmJ��ɮ���%�lwh�#F����p�h�U$;��]X�	�*@3l9t�Cx4O�rx��S8���K�>�J��<�}���T�h;��]i��$7[��6xR��d>�I9�أ��|�`��ʛ�dI�w�q�l��0���R���b3x��g�P%G,�4����
򪄕��|���n9q�Vk���� ���7�y#Uh�[�l� _(a��A@"&wI�ّ���<���݆^ȋ�|�
���9r����vL}d���|���f��E��4�͜��M�J�,7mY#�S�������}z����5�`w��%Gd@�Q��k:h�K����7V����X㽥t�R^E�H0WT1����%��oX,���̇��^�����|�>���'?��_=��OVD�LvsV��PUN��G��e�R�}���W�/��h�/�~�G~�_�������;�X�;���3�m��6��=��ꔲCFi~�q<����`����@�J*�//�P������ٕMD����A{Y䄞��BS�T�D>$!��z<����P�GfpԈQu�H��Q�$�{#�J%nwR����p��X�����8�jcD��b���EhV3�
V��b��<"c�V���a�~V�y��bC�PS� ��1!��+�$kg��"�H�֙N �-%EV�M��^&bj� �A���Ԫ<�;B5�C��w�y�B��b���`��G!^��Z�9���`��p=g�R��y'�1�;���8����֕�,c/�c�����E�в��h�Y�Y�6ۮ����^ﺳl_�'����w�ޫ@KVϙ�����(@��Z9�}\�tQ""H��Y��yE#�lA�|NM��{��_���G���ż���Ǥ�l^���~r���}T��3�z�I*@��z���i"�o?����~
Q���(o������������7X~���Cz�3@z�[�ۺ���"Az�n��9�i�X3Ju\��5tYÚF1�(�F3�(A��Ņ�[�
�yq�8�Q��c�R蚌�AK<�����������XR0/�/?��#O\�0B��_�`:.��A��S5����٘b�b����x.�`��L�������"z`6�S��E9�V��G$�;R�;K@KsSD �i�B�*�̸�|�3�%b�f'���#�a���X�q�Lmq՘�^Exn�a���F.��%���<�������E 20M.U��C�"!�:ӄ��3Z��G#��	����5�bp�d�̀������%��w
Y&��U�̫hř���p���b�m汲r	�d H�)��"лh�EK��;V�hh�n�W�@z�Bq��}���O����%C����>�Cϣa��U�ߗ�S[�P�Mg����>�3;~x���)}}��4M勛��:��oĢ��TTsT�&� 7I�a�u#�#���6:ؙ�?��Qlh���NWۜq�+7�ɾ� _��x6�FD�
��C�~�k��P�^@Q��H� �R��VdңA)�5�ʺ�� �g{]Qfy�Q�A26X�TK���4E��*�#���(�a�,�;b�h�5Ē
�x���49dO��Z96��(���V��d&H
Q(�eR��l@+�iRђ�!���c��LP�j6p��z�M�ɂ��Q�4&�=�FQz�
$2���L������'�K�(�
pGCO"b���0��vxQAZZ���Ӿ���������m���V��6��H+E�݀�6M|f�/-T1v���3�REK�Q�BJmA��--|��}�?�i�zd��}}�_�(��u��_|ෝ��{,QTC��Pw^٪2R#��*"(q�?¿������c�����[?�����g^�����5q(�yec��V��� �;�´u�D)|I����(���R�[�F���A�A�,P69��j���D� �B���=�ii�<�~���U�����%b^ѽ�D�F:���<�R	����ј�=��~ⱕu<���sC]�F#�Гe�6똩WP+�����D���e�b#	���+eC�L~̜UC�K<�$[I�6��+�	���#D�UvN�Pic27P�k*�i��=_��L 5�h	h��9"e@;��3�hs�m�� ���U1�<k��m�Ij�N�>�J�e!Z�.3�ɤ!b��R�Q��-UӲ�Z�N�PA��@,,�I	dv-1u	h%�Z�^�U(8"�1�=�h� S�hi�t���u��k7В3Ԃ�b.�|����?�uၪ@�����e�`|흪�G����-����.���l��qg�b�Yu�z���G��ZQ������q>����w����/�{���(��O�ޱe�E��z�v��k� �@"(�)ВD���d8��g�_�v�t�"G�Q�(��Bհ�jcym�
��Uf���Q��d�߂�(%c���,n.i8^�awm��$�^�ۜ�ޤQ�$�"!�,���4��N_�p'׶0�M��9�������<���..�@��1�X���7`�VA��hBM��,�,"2��$��]v"���N��tج>˗�Zxr�G$!Qb2�hEj'�$~N�v���� �����:�~��E�A	%��*˓��!�\i^M�Z�.��<K�n��sf>ˆMR��v�Q/%V�7؈�9��JA*!�s<o'+�h�H�b��K�5-�Ω�����$��?F��C�S�}�A�1��ץ�K0�hg��w�+���C���U�{��+g`t�dc�+_����g~>���=�J�4�桘&��cH�:��E�w�I���D���S�������w������^�����"�����͝v��Q*�P*�\�R�ءְUb���F��'�\��� � C�5��-�0t�;��� �9�ݒ|����>;?	nM9���{��〖`6r�l���    IDAT� �w�R��jp\�z���j�=�a��E+�>z�4����HVZ��{*˺�b���JSQ����q��[�y�k�h ��1���dC4A�c"��-��(Y96��d
F���b)��&��+Fb���������"i�I��t�h/`%��K�Nc�������\���9�5ͅr���O6�.\\�����qΣ�r"�\�D<�����v� �湗�׸���[�nUзĢ�9� r͚y��b�΋2��{���iFK�*ZZ�($���ț23�?D�S�����i	�j���_������[:�tc#w���u��~�_[�S#�����0[�P�a��G��!����\�G�Q;xx�o��O����y�g�����ҋ����,o�o��t~%�����Uv�d���݆
HEO<}[��=eM�D�������-��<�\R� ;�-��Y-ES�q�����e�
>���P� ���8�b��Hc���w�wt�;~��7[��ŋ�@a~�uᩮ�#v�V�,a!���`ͪ`sc�U���G0LM8�
Y���PLf������wL�����e^Zj��R�N@�iY>��� -�=s�8� \! ��'-�oF@R��0�(S��vV�1W/��\�=��/���*��{T��J��gN3�x��(�KW�H�C�K��1y��N�!#��fj�B*�ϱ��
1������Ą-1��c}�-����:F#'3���r��F9S��s��"ǳjb\W�
W�S�mh���_�ݽ��U{�{yv����W�;�Ľ��X5�o��ZW	���n7$����x�i>��">���죏�����_���w��[n�e��ٻ�g}����~�P�������/Lg��HF	�DD��+�X��s��jX�%"�e\_]߆���,!�/��1�
���ᖚ��Z��7�1�@���{��1�:�B55���f�0M��2δ�xxyOln3ȎJ���t}���(W�(T�x�������1F�sf#s����J�M�������-����8k�F^�+BҠREK�o4 7@ȿ���<�x���3���vB�"e+A��P�HF$�$΀%K��ٵ�HBh#u��ASE��d_�R�dm����Ç9(���u�ә䠏Aw��ůM�J��|������L֒*x��1yl�e�BȲu�6%C]��3��+����Ԥ5�\����JN!S�LI6K/M����-�p�|�+ڔb�"�L	����`�T0k$_>VS�������{:�W��뻺?��9��W��}���*�{�5IB�l�(��|=s&bM�Z�Z�_�{o77;��?��_�?vl��]}�s/����v��<��#���6E�a
/0�#�ӗ6��=���>�H(��v����qa(:�p�^Ƣ�h���Z�,�` ������p4`G"f�f,��G)�H7�������*N�{ku����9Y�"�77˦0JX�1N�8���>�j�V� ) ҋ�je�B�!	��Ok9.N #e��#�iFK~����3�L2B@K��Zr΢j�ـ�l!J�$ �x2��o#��hAf/_�f�$�)W��IU�()W*Y"9�y���P5$Q��C�lX��m��n�S��㐈�؇jV�]��@K��k�w�U������b~�0��+?�X:�� ��_�4�/X:��A>'�Z�`s��@�3���n�k���/����;wcz5����{���<��eI~��ʊ)�!�uN� �8����Á����Non}�m�y�?<�=�� ���X��񥝁�^o��sz�z/���+� ��R�-��^"�Թu\��wr�Ur�i)��P�G�^YF0��i�'6ji7�4�ڬ���m�;��A��"=�Ke*U�+en}&Q�V����3�1�l����P(.NW���+Z��,��g�}�q��c(h�"��<<�Hu��Xp�)I1XC��.�67i�Y̉3T!�!����2�R��x�CƩ���@������gZbP;4Dv-�*�8@8�"qG �(p���3A1,x~�R�ɭ�|>�Ĩ�Ȇ�:L�"I���JAM������������B��ZZP��8f:ִ�e��������gq~z���v��Z�f@+�r��D*�ˈc��P3sM,_ހ���U�-�v�R1������7��!���W�|�W�ѽ̻�<�p����}a<�ɍ�%1��[�]�D� ��d�T��'/_>�>������������˼�{O�
8����������a)�Փ��>� A��x��
�/d�l@�E��Qg��NCl,V*��ܱh��:��!
��A⠅t�G�(��0
E�0X��:���^ce�����8�c+כ�!�+��*�hj��Z��Q tS[���\@/R M�W"gy��D��$DUg�)�	�q>}(�F"�ȬK�ky��,مM�ejA�D���Z���uLmeY㊖�G�Z1���!�>��/�&�AV�1D���(Y*&��&��=!&���y|��q�S����5imXe�Hj��h�n���\ZZt\���V+Z���v����������jK,m�ZǤæ�� 3�xv����\��`�JT*�Rڲf��=�}ܥ^����NYk_={��SO�����=Z�pl	P�T���-r.��p��'nCWz�z�����l��o{B���^�ǹ�k/��u��Ѩ�����}?�m$),�p|ZO�Y�ZkOP9��|)��"��*��An]�Ǒ�����<聏��o{`)"�R�T�u���蹙��Fk����M\��Ѣ�;#�ZG۱��>�8�ױ!)�u�C���hb$0��5$���o�L��Xe9�"�o�������"�lL?�$��leJ��d���jR�N-	��4�h	�	�"�73�=	�.�&���Y�Qni)� >mw$���ca�A�zcT���e&�����J-$�q"��O�,�@<��R��X`g(�˚�<UŚ�3v>t�m�e�r :i�^оP����v�b�pj>�����Haq��̉����)-1�	h��(�hmC8�4~��ż��Ǥ�?0�ԃ��\wc��E�=<��BQ�0M�l����#�e5gl���8���)�����w|R(�z��3��=�ն3?�~l����G8|В���0�7|��.m�*��;�r���)�y{�J�[gjX2%�g�ȶ{d�l� t�s��A��2Zc� ag4���ά��|���0�T*����fH2�by#��zT���=_��U1�Jy�r�Zd�����$2���uʉU4N���Vf���&���(���%��Ky�CJ"�@�
�^,ІQf^A�_��*I���CF,EQ(�"���lu�ȗ��ZEN���jR�[�����xL�; C��i�L�oE��d�@n��f�m�o7оPEK�R�@j:���q͜��2��F#�T��8*�wl���L������H��	�� -����ౚ��w߶��:~��&�����U�>w�����������~��
$Iw�(�9tC,?�;m���G��۪�����_�����O������cύ��z�/��P��P�("$�u}�ϲ�]���v�絊�㶫��Q",H>f�(!��iwᯯAKc֓�}b%�VS�����I%V�/
X����D��V�7[l��OR�V���U�L7�/�у��#p`��	yؒ�u�i*�?���H꒐;�ٰ��*�BВ�����%�1�E�m�R��#w�Nl��F%'�J���h���%h��1|*�,G"B�J�h0�ـ��b��p%Naj��ř�F��b�/�x_���i!�mZ��# �*������T"ve��-4X�3��#�c�h3�0�޼������m@�{NKϙ�,e��)В��c�Q.�طo+��p|�h�J�SK����1h�������~b��+^�7�o�a�kk��_��{֞y���X���`����.����ի�5f��pU3�ox�ZZ�7sǎR��i};�c�9^�g`�ݞ��?�#�0G���^��	^�v�a��Kk-\��"�����F-�qR��pH
� x�v`�/#G���1fs�c��Ø,�Z�ۜG:����x8�n������������
L���]�o��\Z���\'�!6*��:�)e��Uf�Pط��1�	Af�Oֈ�)�RP4&t�͙f�4����M3�hď�\Z�̼s�8�����=�
��"9hn����,rf/�P�L-٘�=�*�9n�R˗&"g�q���d�0�m��/`k{��x/^^��c�a�*�b^��qd_!
=��$���R�U��r��w����|��.X�<�ϖ$�!�.�u�HtuF�;Mg�����~"�B�c�TM���O��E�t� .�вt���*I8���U>r��9{� �Zl)ܾ'����c���"z�д~���}ah_���W�^������ڧ?��;�O�HSUg+i����4��ˁJ�DU��z������s�����r�����yE��N|������C����D�p� ���hP֐j:�Q;N�Q����Z;Da���Bwq '�XD���߆J�q���@$K@d�Z�f��f��(x.�����N��8��"48���fr2�"�
Ef���D�Fρ��2������%x������T1�Qۘ�LԎ$`!2����$\]'�Zbh�H�U�����B@?Z��I�7":eV�4��n�@z�I��*�g$���:v6V�8����8�����yLRN~����`���F����N �<�P$0'=�,�q�é�rZBY���e������U`�*u^\������Ͻ)T�_���5���sl�J��;كv�𳵠�ҧ�N���Q��;@�q`iC�����  (T�S�{�Z\��Z*�����J��Z��xc�u�m����0�9�_~��֞8�+����sAP�� �D�VY�Q{*Ȫ��)(cY\k�z���~׿S�Ξ��k�P���>��c9��,l��'�����*�3k:i��`���g/����@�"�Ʉ�j��tQ�;(��uԅ�� �9F�E����EeM�n����>�V��0��v\<v�"�I���$����d�F��h,]G���h4�j�J��-'Hr�SJ��:�R��N�a_j��b�S�m�Ā�dnOBe�=2����Z����t�7�O1U�����OAW��W�l�BCJ +�ĆX�1�6����d�=��ȕ.U�*�iE�`��Ɂk�7���!��lB��*��"��rb9��L��y�	�u��k���,c�=�%/3вDj�׷����� ]sL�aȀ.�)h�7?�sW�wc���2E%��)ꖌ*����%�˷-~��F��Ca�b>c��Ǽ���+���{��^��\?��{���/E��-eQ��QFT!A�Yȃ�t2%}�t�����_.�[��[o�����B������+�g`yǞ��w~���_���J���D��8��m�q��E��]X�0�I��^@��
�A���c`<�LLWrOJ�)3Fނ�&<���I�?@�q�?s-��S��p�Ɗ��( ���l+�B���ȵ���7��B�ل���	:D��sv�Ë�,� M�*���)�$y�|4j��h*y�J05�Q���D�2mR�%���}Q@�f�$��d��Խ��^�r��*-g��m���8uV7����[�D$�Hdb�r���$U�-��΍Y��)-t���g��@+R���횊6z2/��}�@K�rR �|�ԭ|̕Xڇ'�:��+�ZD,*� �c����K1����͕��M��W�T��{^�{�k�9)���у+�>�s�K�ޟ�D�G<���V�?|�ʣ�9���4g&��k��|�7��ﱴt��ޓ��v.���Q}��h�E���1M7D	����L˃�������($!�r�r�#�n#�nCt�=R�|���7ᎉZ�c�\�&���N�0����{=�o��)*�� g PU�)9F���J0u�Bc��0ru<�҆�8��l V���/2 ��D=�����e�|��2�d@{Hx���b�UYa&0���ΈA�3]�����5���ҕ"%YE+�TaҖ��\�+���w�#v�BpP{��@�ׁF�dI�ih��� ���@m� �Z�MɅ����WL6��z��Yhy?���@v
»��g�����Q�����6в�J�`w:Ԅ�pB0�|���ǎ���}��#�J �)��5ڦ��*z��:����;�w�H�ӧ��s�ꩧ��SO��EU�9*ͥ����:cD8Q��5��9H���凌���g��[��Rg���xþ/����;��}���7�n 6qňi���CN��nlB�G0�1��E�ۂ쌐�C6B�v� K�T�"#Oz��~"���Gc�0����.��Hry��X�Z��㺰JeT����f������9������XB�V���P���کr�٠b"L���pv��*���@��%����ƚ�@Qe6����L4�o)�� V"c&
�p����6�hS[�,IV��nma4��l���V)�w=�\��������g��͡ 4�&0M"L���SE�^�z1��e��k	L��)8�/��sIp^�c��+k��BSbȱ��Z�?�/��(<(d��6NBXZ�������a��H���/�~�p���=��������Vþ���<������,{��F!tJ�PP<{"+R�XzA33G7�a��P�#�t�m_��a�y�����q7��u��A;�����e]�p)���e���n����ڀf��^B��tІ�I�#�U��CL&I�Փ�]�Uآ�K�>ζZX폱m����	"E�K٧�ڮ�Rs�����&f�M��h��;���P�w-_�+��9�Z�NQI䤈����Q*p>�TƲ�e�$�I�G�[b��ܔ��	TUE�ʞ۸�W����;W��0ܺ
��:�ߋI. %W+Z�R���9P$U��n'c+
W�ł�6�F���vs�Qh̢;r9؞��+�$�@�崘 �i�ɸ�:�����k���^�@K��-��UlI�
+&�_�SO��8�@��1%YZf�XӁ�!�"�_�m��[G*Շ����z�|�M,d\�0�][y�ٯ=���V�6��&��e�a�*���M�np��Co�1֔�XNU��co��~�4����� L�/b���=[[�F{��7��W��S��^sak4@���h�lG�Z�0����F�� ę8��SM�UD��E-��#J�*c�q���6.t:x�4�����*/IE�Z�D0J@�Q�ԀDD�1���~;T����ÈsZ�DY�*��(�@�S!aob��~dw�$(b�˖�٬���d���B��]Sh���ٳQ�_L�R�}�e�*�`x�N����5&��P�E)�.͡�"b�E�Q-er� �^��Ǯǖ�� A���!g�y
�\%<��D49V.�w��CR3�Q�������3Q|�W��>k�κi?�yQ(�f�*f���Fω���`�J��4�j��K4��­�J��P������{�zսzz�]ܷ���m�=�����1�Q�D��>4j�y.��Br)J�#[���?�ֻ�C��g�M��:�3�������� ��	�(ɒ�؎Gq��e�*eOM&3��'.�T�ʟ�o�������k;��N\�d-&e��L�$b_@�����}I=� )R�ĝ�[��@��s��|��>���%kjqSYدn?t����vw������{ؒj4E9M�]��dk��md�!�^]KE%�aEM���,U�1��\͐�1݈��C�I�[[�ȶ(��q�LZ�����m�4���T��Tk���$m&1���B|��KH-��u�XTS��(@�0��M�ȋSL��- ��\Vk)�Y\�8��EʖqQ�o<VG��L��գi�6F�~���zYI���`1��z��b    IDATdT�G�UL��QOl�d��wz�Ͱ��&v��X\Z��^M�ݷ��R�E��H��V
�-���k�z&��L��z��u�7�}�g�GȈAE�aj��i��L���C˸z�&��� �b�0�	m$�)�)��V�z�@����Z/�W���}~���v�ko�ؽp�7.����7F^�
��ӥ2��>�.�r�G0�����xϋڨU.��y����=<}�'��D����~�O��ՙ<}�H��У�x<h��-�n�@��E��B��ٚ#��zC�,B�\��3BZ2��f�
/�Ћct��~���.V�:���a}��z�M�'6{�6+Ն$��/� L����,����&bg
�Y���L��IL���� `I���Z��lV�œ�՜R�T*rV��&P$�7��=mIO� ��8Na:q_E;цN�i������Q�DG+`˨=��f�:fQLI�7� ��
ʦ%�T�~����5�`�m�
L��J��v�f�����www��Es
ʢ�loczn���{m�?��L�a��k[�E�x2Ý����z������eׂZ�h2�}��zݓ��-*��w��J3dI�b�ێ��@����i��x� E����ad�8C�V0WV0�y]��:6e��O�:��a�����߽8����K���@��kwΝ?v�ܹځF��;�����eW�P�T��t�ɠ՚#���Q�=�.,���S'�Xs+����`�8����y(�������۾~��hk�Ї6B��{d��bR�Ro����S-ii�*#�Rq��r����ּ 7{\���Z��v�bDܳ���0|�8��pa~E"�h��J���p�[<4j�B2D�JA~KV$L�`;	�E�2�,ޱ1k����k�M[Ɩ&LcN%	��\'@+ٵY&,a� ����=�q5yhuq�"���z���:h6�p[�k�y�2o�V��z����5TMhd�g*J�)	��T���Ѣ���^�LOf�&����K�2i��0���ϒ��\E���������AZ�6� ��Y8���Xh��8;��0�f��<S�Pd�;Z���c�n`�b��|���)��?����*��Ǫ�{�y~�oU\z����������~�yl޼%1dY��WIQ���kVD���Xѐ:��\o5��ZeUk4��.N}��#_��ֶr�P�{��/�#��-�W�?ݾv�WGk7:�n�������H�!�q{��Sٜq��Y���Tk����H\�8�����C���uz����6��)��8���*3_����98nI�0y�m�ZA���"��Ь#�q^b��fb��y+-	I����%��U��V0@@��6� ��-�E˘@K�$�y��`VyqF|��x��z���S*7n'����ض��7�$�C&ٰ�aQ�'�����m#�t������Wp��	̯�0ds�\�8�E���r��R�,,kF�ku���k�cM����mz/�a�v!�hy~�V�o�i��-;A��#F�XjU�0?��0���z���m�4����rr�4]̻ZR�Gs|���=���~�x����@���S���>��G�yby��n�?WMF#=�%��3[�����2T�=��r�P
��:MJ�y��n�W�+���/.?��ܱ�n��;�ɓ��?�z��0_]�Q5�ן{��έ������d��^��Zl���9��)�	C�a�����[B�iP->XѲm\�n��՛kX����� ;q�A����Q�������t-���Y$�ݪ"Sl�m�:���~�ܝBZ�FbOI5�X�%��D �l��<Ԁ��˙أ�H��T�B�"��0���X�C��E�$���"��O�Ο�>9�%1$^����PQ���YIqC��=�%�p �)�Y�d���b��9мbz}��0�q��-T�05��0J��> ���sGf��s�bUI�Y�Q�H{���+W��\o5���l�Z�����ZyoJ�*��h5�yP����c�e�%,�Mc}k��!�܅b�C���b���U���0z�9�~������[0����#曛��}�K��������?�c?�05U�u���-���0�N��N���ΐ�DU��@��aTK�!VT�)��hg�8�թ����cz��8��0��{�yFo��}����� ~�ɒ5ϟ�����׃Ĩ��jYX�X����ci���e)�B/Ja7������Y��� g/]���6|>�tf�"F��֧�k,;���h.6�>��@���Ԭ��j"6ˈ�
���(!'���=��Є�#� -M��g-�9nQ��e9�-u�]�lCRt�>��tjS%���ۊt&Oe�ȏ+f����7Z�.�J����@#8��&��6F{�H�E���VrP�����斏Bq�0Ka"S3k3/	��z��]LO�²]�Q$�;����1
|�;��? �4���8=3��ұ��t,���6C�0 �i��|��w�¾���TL�ʹ���2TbTE�F�˲��n���s,�����W����O\zqh?h+ڇ��l\�4�'���|a�����}�С�V5��D�����F����`�)lVi*�[�9���?�\'!]W�r�����M�ٸܜ]x���z�:5�a/�������M~���ܹr��;�y��Jgc�g�?��щQ{�娊��!r߇�db�H�+�RA�X9��i*4�DfҞ�\�u�0-�F16n��`{�����hP�%�*��4a�+&D^.�LT�fEZũ�@f�dj���4�f#P-�ZIHW��e�6����e��ak�nH|\E��iU!y�M�8;q��E+N���@K�V�#2�ن�6�d�f2��V
؎~��>y��!`s�Mɧ1d>B4�!�8s���8�s�o㡏}�fI�,�L�I���o^����&�i�6�A�r��n�ʵؑ �����*U��
�Q��e�)U��.��>�^|�!�k/�zEKg,��م��BI��-@��]�{���Č�����nƘ�3,�M�����R��?3���ܜ2z?���S�{�g��x�[g�>�����-W~���<��a���82��~k����fOc�����8��*��~�s�3�f��*i�j�T����u˙�9S_Z�jmy�Ui�?��(�O~w���|T�.�)��������l�C}�r�|^�Šߗ�F�y^�~0ܜ3���#6[�$iR�et#�htgRЇ���cc���nW�����c�R��ˮ�"�[tK*W2�MS��<ѧ2]%��U��<��6`s�A-5�(h�L؄b�b�!>�IM%Hє\в]+�7�D9���]��ŬJ���@��m�1aʛ,�h��I7%�H��l���X1N���
h	Z�:BT&_���4T��i���TlU����.f舥[8���a� 5˨N���a���\�s��%o�E2�i2B[LMC�Ւ{��9Þ����@!q��:�->�@�&
@kJ ���0�@�vv���;[���:�N2��M+�B��RI��I��Y�����Z|騢����������Y��\�旿������?�ڟ���;priњrm$��ﬣF�������p㘭��R��t��s;��Ao�ƝPS�����|��ɣg+���j�Յ���G?��{y�����[������WN?a��g�0=�{���3g��(F�(Q˚g>R�X���RQ��NS3�i�g���v�^�5q�����׶���`�߇清��$�TQ�*
 mX�tSb�b���`�ڨ.���V�8��$М�]L���x��X Z�D$/
�lBv�8v2����9+���V'����z8/.�b�K���5���G)k�l��̂�f���P�*�Lo6����$Ce��?sx�,E�Ŧ�z�r/]���0��"'S%0(ؾs����ʊ��{�!,�	�i*s��h�ZE�Ӄ���tIܣl�ǰ�eO:o�u<a;�J�5F�N��=��&��\5q����na���V�M5���搛# ��ru��Ut�>��� ��T�}�J,���u��敒��[�����/�tRQ>�\�}�}/W��s�y�����'�����_l]��3�,���O��u|q���~��6[�b OB}X�(�+ˊ�l�TB������!�R-����v�O�M�^��Wk���oή<�Qm裪�������O�6PA���q�n�M�l�>1l��k�w����$�����ZJ��Q����k���V�5�2�bk�-���|��26�=$������$���&v��n����.�#���E'0e�9%�XW9I-*C����.����j!1�0+�j��x)FIQ�
�G%CY�k>��Z�x��u���6�]Uh�/�Oc���ٴ��M�3��QuqA�H�J�<D�P&��t䯋��B���a�����v_���B;�>ɤ�'�Q�ؗ �agW/���a�M]6?�q��&x�c��o�N_�ˆaa8�cqvZ�:�Y�޼�f�&�&��i&^�{ݎ��oon�ҜF�[�F�"��_ߓ�F"lmλ�J�3�J'�A�$*�
�sc��49[���������s��z�tn:LѨ���y �a��u�fU��4]A�V�rԵ�5�C��ӟyp�_|t��P��z�����tB��֜�{����G�?��я�ڻ�7?��?7��m��B����7�(����FE�HXYx���Y�O�x���@7/I�T掻���u�5uè�_0��E�Q�^~��.\w��y���Ő��9�J�u��Y�5�qm�����F��?��I�j��nIg��2�BL�Z�SWY0q�23b�F��	L'9fF$1�R����K7n�z���r��[���"O�ٟi*�7�f�ck�y&l[�	��3�^��L!�����Z\�9�SyL�	�b&�!mL�T�j��_	��W�j6�b[.
P�uH�m��KG�t�f,Vy����]>�o�c����"�bo�@Mǯ�skqoRE!l0n�JZZĄ��p��u��=,<"	E~�boI�-�^��Ԥ��c�ajd#�@��G�	��
�Ĉ!�,@)���I'��Z�S9�\HD���}1�n@�~,cr�0P"Π���o!��ǩ�Q.YX��E/��O1[a��dS�h�j#tן�쉹��£K/*��s���q���scc���?����.�O/��§�4�;�r�zhe\F�2�zCD���=�U�ľ�,�Ʊ����cEC;G���8�NV�w��c"Q�$T�(Q��b�m�q�f�v����l�OM�]�����Rs�Je�#G���E�F������]�7��A�_��nτ;�۩r�wg�X��w�γ��f8z�9Z�
����O�v��PƱfl/@� �U*#�=7?��Z�m��RA'�PmM#��l����+�7p�;DD-'E+�C$�r)�-��ecŹ`�kR�xdF�]OjV��=?G�c�hMD6!G���{ �I�����-����	��r&Cy�R�R63�\��4��0� �{=�L%-G0�H��g�r]��{w3�y�X^2,A*�4A�6���D�!a�[C$�!;�/����\�%��F��@��ZV���V}g&�^����m�qx��w��߹O�#�dۤ�aGf�wV�k��91(y�Ջ��8�yt�2	� �J�꡻��>оs�e�����yn��?��|����:���n\�����O�:��R	?��O����na��dЃ��iMC1�D)L	L�7��OJ�-�PC�Q�V+�:M+���őg8n�*��5�]7JΖU�\t�sW�z�7;w�;��R[�1;(���$��y���;w,��]�^T������iu������=�x�doN���+e'�ŨC�d��l�Q��q6Wp�,�n�V$�:�$��X�qi*z���0��+�[Sh.-��������o��3��`��PlG@���n���Ki+4搲E�2���*�-JKHO�b�Xs�P���`��(z� ?��О�&���Ū�޵b����@�N���h' \X(�3@[����=㊱�Hd%��B	#k���Y����KS0�����k�3S%K*\����bi�0vz#��'�$FQ�N�C�$���E�~�}�:L5��n��D�?�٠�E�^Eo����a��]B�;����8Q~4�h�5�V���>|���[���=��\�L�iw�1Ө�����WA���/�:���{RsuI�i������o��r����:y��_��t�����Yg����~���/_9����ԑ�x���6�;�mo���bУ��TUjD�'D�$lK���	A�TULLᒑKe���8K�(M� I�0�G�e�L���������A��z��iVj[P�a����R 3���}�'>ps��p玍8���9��p䙣^�6�gS?�(Yr�������7�Ւt�T���(%3�m��X!�1�q�$���=�P~�ϫrc�[i�(F?�Ӳ�ZC'�َ�~���/,b7Ipk{�_~/�|Wo��$�r�b��B7��MP��I�T.F�jBъ�|�QBf���硸-d�1��r+��T�G�+�S���T1E�� mQ����ڻnI��8L����`�m�J�ې֭&4��7�k8��H�Įe �aw�:�����CϹa�p��m�>���^�c��C�h�"5�N�������Uq�v;�7[��ŭ �G���F8���e�RNm�f#R-$�8)�@�!zGf�o�м�@ˊV�	������_z���|���3�'�(�q�d�0�ɛ�U̕�!�w���3���:����G�`���'G���ӿ2�agg����z#�pba�~�8;x L5�4u�;;�;mq��\��@�U�=�����b����p�JBB��Ȣƪ��Z��9�zL+R;��t��g�K}h� W��[�t܊{Y��k��̶^q�*F}�լ�ʭر�%����)��R<�x�N΀EZs䈁 ���'U������E^%������l�s�?���^3���h�̢��gi���v<�IX�}�cQN+D�M�\d)� �ju�=J'j<m�B��w��H�h��-�'i�Z�j4]��j;��s����� ,�7oa���׾�μzN��u�,�^��h�z��Q0*\���VC��I���3n�hra��\�Fzuzy�� �
� �n��@�9�:2������"m�*ډ�aq���@;����moul�HR�:.X��'sC�Y�C=m0���z�mm�Ys1�q��C�r���`}k��99q��K�(�}c�n���f�,@+������i�J��~(��P1��W�Qlf����a!��������F3���u�-7�n I#,�4�۽�/�ܧ����߽$3Z_q���l-5���c���Νo|����ޟѾ}��������_����'��v��~ޱ��nw���n%�6�m�:q?���q`f
S��;�.@�"غ�A�[T��l����̏bt��T�8�LN�Ŝfﴢ#�$:QI�� ��zs
)]˃8��$	5MTM����;F��s˵��{�i��9�mw]�-/״T��@WM�(�C�q]�SӲ�"g��C
��6��	$�+y����$y�皒ed��A�XZ��0-YV�;�x�Q>��QQ9��f�y�Z�Y�[�s3��
{�
2GRO��:	{�D2�Ϩ�Q(��8�q
�K��%����騙�0h�`f��A����vs���J�^���f9�KOĆ�V�"RU�|���x敳"/ato8������:L	��˓!6~lS�YV���H]"���ܮè�Cu��u�paUZ2^�9$�diȔ h)���7Z^�w�o�rǱ7���:~�,�~V���[ǻ3JɃ-�1H>+�٢}O��#�3��)ﱵv��e��l޼�<�0?;���eI.���_� �RC�5#W	�w�naws�a��5	�`W�s�N��A�0���P��9Z�iD��D1�1�4��&����ay��4~#�������}�+�C��)���;    IDAT�;6�ɓGP�8��WΡ���*�J��.�څ��Ū=@���?zt�w����*/d��N_}o���<W^�|y�?�����W���-M�D<���AgG���8�����C+p��OD#_�ZΓı'�D�G6&gz\�=(S�ql��Of���\as7�-�xÅ�m�"k��*l�%�*S�W3��<
�$L2NǴ���I����鱦�n����1���fj��%ۧ�#�2[�1R [Q��J�{�ϒ�ΒL�UU���QS�T5�Y��J���<�F�@n�yf	;�4%M�<IV�B�h��m�,O�$)��c���{.	�V��" ��m[&t�"-K!%ьA��If��(Nnح֥��O:z�y`�W��i�[��/���<��g�����:T��\W�%��@Idk����v�pݲ$0Gְ��^�ds�ǖ�V�;��'�U��]��\�a��OT1��ٮN'�y�����c�0��;��� ���@{?����6SIS���ϒ� `������ ܢQz��t�FY�{[8�E�:u
q�`���C�|� �p��y?� j����/^8�GzP�i!�jt����&��5��s�t��WPiΠ>{ �UE�2 �I�l�>�8�# �YLr^�Z���cڪ�82ߔ���7ױ��0���{���\�����Y[��;���#���rj��}y����?����7�y�q���C_����s���g��;���5)S`[�ڽ���J��cG�ⱓ��u8���#�W��U�"d~(-+�Ϊ�ߕVh�Q!40[��l��,�e�t/�fċ>�Dֿ�P�`:�T���F�u�0�\ղ4�2Ӵs�~�*W��~���v3M�4�̱l�4�<O�<ϲ��|]Qr&��Iu��M�XN�u��L�gqƩ�G���J����b'���X���2��A rz�r�g�/��ŢI�*�U�䊃=�s��$^�&��� �7�$�:������N|�ģ��ò�n�j�������}��g�������/ܸ	�4a8.�(��-]��D��	4���[0�
�;)�ܖ�
)��,���kP-��m�m��&-eմ�)�=�m�-q:Hi�T���lSHC� Ȩ� 7@ȿԸ��t��؉v�����ϼ0�{m���-�Q)�"�)�(b�P���/t���M���#6��T�q^��	В�]j�҉ �^f��!Ֆ��P�s�����5�޹��Ǐ�G�-t!��|����g������9����L����مPM������hi777����jk�)��+boI�e�����,)Z�����<| �ͳV�uD¨�t�0?UE0��b��C������R.�B�T:$C�Ut,������Ɠ�k����_�w��@������j?�쳳�}빏_�|���$��a�[��c�J�=!P/W����x��A,�Lc�ZA˱�z��e�!���صuMX�l�E
%� (�@���e���Q�!!G�0B�̗�E��4Ŝ=K�Mk
CS"�teE�o�ʠ�fH PӔ��b[϶-$I�((L9��;�}!ט�WE��,�cG ?K��	����%�����}ƪ����� �.�i2�%hKE�ih�Ρ;�0��<U�$ӵ�FY���y볇�X��9���|�����JdF��VI	V�Ϳ��>�_��t��#��:�f�$��A<���dӔ����4�q]�����aP�cK���-�th�i��Y�#`�s�$.O&��t�p�Rδ��A��$�]X�j1�}��6#��@+�)\l醥���	�N���,v���?�o����X.ʱ�0�a��"�F� �*z���)Q�We�i��g�Qo�p��u�{�*�Y�x�a�W��HR�w������i�1����s4�%�j��ќBkvC~���{�C˶�.�r�C��k���5n�:��y�����麋<����,�[�ן~AX�^�"֋�g��6��k����<�������Ϲ�H��ӧOO}�_]9s�����sa�A���ʬ�݆k�����2�X\�g?��e�LuC�M۹^�`���ToB�a��>)Z��g�?[���(Eڴ�c+��d��������t��*AߌL��E�K� ʏ�\���T>�X.#���y���E���hL�!.�����@%�d��_��6�la��=�*��&S�Ug����j׬�;^����v�9u��G��\8��LOwC]WgZ�m4�9L�8���_�������~�?���;��æmY$�M���ka�5�~�sw�ȴ�b�:L��MQ�ak�r�UC�u NeF���Q�Z;		I&<*u.
g�,�Z^Q�ѵ�f!�x�x0	��,G)�Sz��VL67��h3q�z󊖭E�6Prm�&'�в�%�N��4��y��"�����R�&���z���9s�/�h��6T�:;�l܄�z(�@�&1����T��ݾ�8�:V���1�d~���kפmL2��Ύ\�%�B�"�(�ι�Ԛ���{�mV�вkP��q������3�X�\�p�E��hO�,bf����/c�k�h�f���`�Z�̨��O���'�Xze���HB؇�MѶ����?>��<��՛7E��UӘ�<���ڨ�C8�A�`^�(D9VZ��Z827��VSro+��D)e��mIgI��g�&�V������s��*��T�H9ߋX����OP�h�n�=�i��G�kA]��4EɲE�jH�)�"�e������I���Xc�I��2��CQŉ�Iܐ4��:|�6H�)2?��LUc�fCE�.5�A�_U������3�wZs�d`w4͟�������S�<s�?��_��3�?��� ��Ls~䇭��i�g���
�V���i��[�e���R�H!+̄jU॔�Pi,�9���(G��8wkG"�8���%�KI�#aY&L��)Mb����	|��Bz#YR<"����+�	��k��<���Z��PE�$G���i:(hy\l� ;�tL���	h�EG(��Nl"I������l��c���B�㘒+�3����n޺-��'��0�#ɩ刀ٴ�F�%��*-PK��D �`�)�AE7Ĳd�ग़ m�Bܺ;��8��9�@~wӉ�*�-�m�r}i��#�J�,����K2����mǚ%��IE;e��6�Q)�}���3���Oxe����z��^��ϟ�������o�~���^���^���i3i�(�h��m�{Tx�R&y�n�h�j���f`�Y�t��CsӘ�t8�,S58�%R�����"A���,� E��`$�}�M�[�U���@�m���֬�I��(��!��VT���@W��cr�df�������8Z� )e`Wެz����DX��:4=W5-��4R-k�Y� H����;��S�a�g��37�-�7��*�L3F���nh��z��/�����'�޼�p'˵Fc6U�*�Hk���B���k/9���G�B߃�[b,B7!kh�G�a�Z������Q�^D�5é�?���S\����ZZ��I�*�bsc��JR�\��v��,IP�CIӻ��������X�T��qr�����r�伽���w�h���Ɖ�Ǿ�d� �#7V�*#��iy3а�H0���ջt`��A���h�;��ػ�.�2�Y���*�H�"Y�vJ|�I�#��J~mzBX��U" �L���Z�D�eHr��T��m�y-��c��p�ō�M�h�:�TS�V�{�ӎ������k�:����Oxe��Ch�{%ϭg��Og��泏ܸ����`�D���Y�Nš�n�^����T��<��b���\�_ޙZ�4l3���M��NU�4�+D���W�9�r���83X��
�H$���˩�ym�DnF"�	��b����Y�	-�D���<[�$�p�H Og�"�Yf�� ,	KZ��p�;s)A�sa(�Ut3U��<%�<�F��7�[�F�Z�U��;�m�)������^�ia}f��C��zUG�f�ľp�Ճ_��Y��_|�ʕ���q�<
�y�qjI�8V��d��Ŭ���6c�\�~�W� t�l�v�8(�i�ab@����Sb��U�g�`U� �D�?D��cm}�nIM49nl��6�w-T�$�;g��ppS�n-[��q�E�)C�:�l�!Za��:�7��N����P�5�dd >�j�V�?�5Z�#�=��I�1����kM	�	�(�%��̡��KD0B%�5�u1C�i+��p��ښk���#�UzM[HU����
���
�2 �f'�`$��/1y��O>����m	�<y�n��F��Ψ<sT�G_y���?�|fh?���C��vvv*��s��7O]8w�rMy�p��Ѱ2�.�d��'�3Cq�O�m����e(�榦Ъ��t]�J.�4���(Q+J�z+g)tV���bXtA3Z	R}&�hL�:�H�G�iV8�7B�TFo8@���0e��Ĕ�`��p��|i�B�J�,�B���i��y��
͇3U3UU2�qs([���R�^n]ͱ6a���/��j�u�9�ة����{T5�8N�UQ.�8�*��ݭ�7|���o>���g�}����'F#I�0E~�);�r�&V�{�896S�\�zaf���j>Q-W�(�!��#�5�N��"�Mhn��,�+��2J�&Rg:�:��:�>�l�BW,!7� �}�U��Z�	I�A�a���`<��_*c��Uъ�4	h��U�M"OZ�Z��
�v�K1���lK����F3Z��	xe���k�Z)�j��6XM�:�mܹ~	٨��cJ�A�,�$��T�j�p�5I����b��X�T��7l3�pf� ��T�U$�Pb���.F0��ӭ�J�F��h���h���e��1��DH�hu�������~�� k;��c�}U��pmY�P�b���5�}�p�w�_9���?�h�!x��}���3/,�z���]_}4��P�e�Q7|���M�p9��bQ�a�FV���+�$�b���c�����w�3�:��]8&i:�d�)�<@�㲅���e*��%�;�d�ұ���V���������'-f�4�(��,�;��Ւ,�c1Z�O�8��4�e������4�ގ����fl��c��M˴黷
]�������u�v�Ug�T��陙��*���]��N�䥩���tϾtef��Z�+_{�';������Q��V�,˪�aXJ�X/�Mxް�H*��� �H��q�0e!��:���J��#$�&Qb��bz���%�zp���[B3�y�O"ل�"
���c��ưI{_KFnR(�q�F~ �U��ĴEk�@+R,n��@~�ֱ���&c��Ql��H%U)A~��b��J>
=�4jeX�"6�܌��5�f�
��4R��Ռ�H�-��'��b��/��o�+i�h�EwF*�Cqx"��?�a��OC� A���^���>�8�0��(�x��9�a�#G��֚Y�d'�>%S�@ׯ^��ޞ�'�ZSH���x<�(@V\ǋ���HnF����}��{�PM��ϵ�U�ZO�6�d!�t�_��g����̹K�*��D�����a�hZ9�����?�R�����p��^����y�+�ˣ�.>�}_z陹o=���3.}���֧{��IðIT}S
D��P[�2�{]��%?c�WX���#i9�,JxB��
u��m�T����b�1Q���1�h�4�kp��eG�\�1٦�x�	��,D$r�alv[ѵ뚡?7uE�C�P#ðo�J��@���Z�(z�+J�v�p�4ѵ�.�ںYNM]��R)�M3W-KS�K�([��}�Zt�}�G���V_��R]�}m�q����g�.^�r��k��mn���Q��P5��fYUU'��~&3��WZ��[���+s�����}�lN�l��#��l�q�Z8t�N�8��O<!���.3h{�H"!�l�,�g(������n��/��mXMa��.NEbB���ƶ�"++��o����U'.O�?] �u�׉糰�ǳqi���G��t�r,�M#1��-�ԥ�%���&@{;1M����[�Dה�2eM��+r,&��BFir	�TB�S�ť��h7�]��Tp�Ă�,tv�R&a��4�z�<�=tR6�%�&"eS�e�([�j�PR\�r	333���RM��|�8s>BҔ|
v�#�]<a���Ip�0������d���d�0��L�߄|�f^�E�赛��oӍ���i(0���AY��?���+�nbs��Q�c�ϡ8!�h�V����e������?}�~�X��wq�|_zh�����<��K���>����/���o�p�?�U�GL�t,M�F�?�Q�ŉ�0�$.ӌAV��h(�?H��l�E��d�9�\<�.�HB�|Y�hv�E�U�I�"0{�v�ҐD%2i�Y�BԁؕR�T*�P�V��Z��ԧZ;�cv��Hl�̃(RbU��4M�J%L'��k4B�~��O���`v��իz��?���f��1ow:�յ������z����N��N��t����5�8��s�A\H��N��J��8 !^��3fF���NO��
�(�z��X�Ztu��E���"ln�
�xaa	�j���O�9}�YCcf�v����ǹxLM%SSSa�4��$@]歱�0�q�ʪ̵'�	[��# E=��,�%��+"�tU�x��z����7Z�d\9><ۯZbsٶd!f�+�Ѥ�h�z~[@�'�	�o
9Pю�@1�Ȱ��a��؜6���NV,k�e�K�2�$9)��x��tgk�/_��O��D��֜�t��[���
μ��8���SpS�* ��I�p�*n�p�s-�0����=�w���$oh'`�M�k69ŕ$��<>���=�`��ѯ<�W�l������N�Bu�H��.��m�j��o���?��o����+�Ί��?�>о���]{�?�z��+��/��y���mo�}B��c����qRͲ�"��뱐r8�yp,�NY��-�������4S�e����4is��0�{�3��D�F:�������(�ִ(�W��ok�z�v�sn�te~e�v�T�6��r<�lhS5�N����U��4U��_�U��W��N��g����k��X���t���a���^oio0<��t��k�y�a�h������gyn�Aibd��X�5��%3<�����WN��H5;0\�� S���p�E���q��m+���9�c�N�ޚ�'>�cR���T3p��:.��pm3�����<�<��m���S\��*��v���yT�!���}���ԷrF�v����\�I(+���	�e	*��8�iE
CM$=�>�y�Y.����R������+��aڰKe��:�t;�[�����'�M� ���077���:�ʎ��V60'?F��Q��44�M?��)*�6���d|%�Z�������:�j1~�g��/�G�?���h�
�Ra�hk9Zv*��f������o����^���\o�Ks/�>Ӻ~��ɭ��O���Y���ۊ��Ǳ��1���$��*i#P�T�e:�����6�q���0�Q�i����V�!�4�����z�Եtf��ۻ�8L:���-?	��U���f:;5�43�2��ah$=%��$N $�n�KO��YbF�'qu�:T�0,�D���yE�Բ��VƖ��Z��(K�d��*Lg)�x����ݱƳ8St^���X�)��2�����h4DQ4Pu��h�6�S���C�>��C���إ2��T�b�����nq��JE�B֙T�vh�8�[�k�Ib�ar+�oQъ�GHf��-*�	�����[���~EK�-��he(���� Z��Һe�<OW
0����[�tR^�f1Ԝ�����5�!�}-��[�+g_�Fx��_��\<^qb��mtvw����V�&���pkm�zZ��^q1Ӫ��/��v���?�u>��0�M%Y����擯�0��^��~�{/+�7Z�W~��������S�~�.\��^/7h�RM��,-A�Jh+����/�(����|��ZV/�Ϝ=7�~{�����	�𨪨+P�z�ev���    IDATv�fl�b�ܵ	,|����e;tNb�*]�&-*VV�ŊDc<{�{=�]HP��9}��LۊtUF�(�s��F�(j��A\�U�(�8kV2����8�,6�T�4Qt�Т0���H�.�J��F��F�F���R�HIΘ�ѝ�?�Fbb�A�$�M��p17,Z�b�Qr��H��� �k���j�����S�N=}�ȑ�����-���7�R��m�p+�)FQ UY�+�tk�o�����2Z0J�"Ђ#?��ںT۔]Ml{nj�:IȚT��ԀV��$o�X�3�}U����?�,�I8��C�3��M*�
�狗�H�w���T^���2�nm���073�!�y�^�����v�:f��8~�(�76q��:�<r
pje:B�N�L�!�ʵ�p��h�n��l��6�}�Z�o��X��*t�@�d�T"|��#������5�b�>`�jP����iĨ[@�QB����/��������K��:�^?�~���>���r�u�Ν���F}}{{ags����'�$;���AM��q;���6�m>�H�)�	�"W<ԭҷx2C���Pb��Ŀ����+%�Alg�-�d�1KLÈ���4!=�TKMQu� X�q�[�-CM��n��kV�5����I	�=��"�l����T���j�"Qb�f�3V�Y<����"�m�ˑ�����Tk��Ï���O<q���Gw��||�R��Ԩ6G#�������k�����e7���&MB��f/_����C�z,�J���ɬ�Z.I:ڵ��X����@+]��w� [�����J�8���+ڻ��;\��$ �|��PE�����&�
QΏ*��jّ����&��]���ek9M45�d� ՘j�ZkPs3(lz��2��GC̶Z�L�B@��ccwgS4rэj�3��O~�Ԅ��5�YBTLIQ^�������K�����ԏ@�q
7�k w2�8��1���v{bڱ��9j��Ɋ6G�Fhz�_���<�/����/��9��Ξ�]8s���ٙ[��|h�N�����q7�L5�$q4Mc�V*]a'{C�ɒY+Fc #8vz#v�l��F��Wg�w���c�%����
��Q�N��O$$��|�.�J%7�Ɲܗ3�	#���w��Iۛ�yb�A@�����Ŗ2�C���,K=˲=۶w{�������C�+�;~l�ɏ?�}�����������_�X���D3���\o,t:=�hR�*d;I� ��!^���k#�a�C�L�IEKp� ���7�g�J���Ia{m����ԁ��2�N�9&�:�}3w�4�����=б�-L:8EQ���E�����������0�y����Qo %��v��h�G��Ȕy�$������}ܺq}ϗ����}zu~�#3\q�b�?��!�SXA�A+��
hy�#O6�Zsrm�&�� ��	�;� 2>�㇉�N��>�K	ѲR4������Y���}���sϕ�_�V[��3{���ǒ<;���b���$k�i����m���E�F ,f]� � 8U�K��Z 4�'�f׶
;�4�#۹� K[W��H�!���+r��b@��]��TI3*��5��=i�Nl�D�K9�h�q���
���O@���iC�iz���i����8�Q����j��X�T�kO<�ĥ�9���ɓ�'N���m��l�u~s��ȩT�ވF	4�?0���{^���;�xۓ�1���5=i��� ��K�~�,�l�O^�̛�ѕ4%i����Z�bd!���^�D��h����:x�̔�IBQ��#��v���r6[)��y�t{=,-���/b��A��u\�ts�r��;m��.��V����54�Ux����7�u���a�C����i���W/� -���̀܂P��M��:�  --TE"d9�՚SKpdeNZ�[�m�����FaZ�-J{J
*Zg���@����{W���ӧ�;�A�ֵ��+�.��޸yd�Lq8���4���,^D�Vt]��(�UUբ(2t��4M��4#�hlFL��kY-�+�֐�����K��}%��Q�lE��]H�����!Eb�&`JֳH2���b'>v���Q�W�0d�]����I)�{/��=��n:�{�Q�]������x`��Cwz������C�ou�<�6�������ޯDY^�s[�I����N�#B�X�7_���7��;���	p�Űv��shb��flml���d���.:iٸ R�2�8L���@4������_�_��%@�D�3Fc�߻��t�W�b��Z�rD��`Wy�[2��{(�2�ڔ�ou����~yɽ�������'/������̑�ו�y6���P��\w�g�K"E'�)��b�;�11;�����Zi4�IdW�hGڡ�Ј��DӾ�ڔG�`H��l���$�U��.6����������y��sω�{	��r-��
����.� �%�܊R��f�3T�S1oj�on���<Bo��nP�biiiI~��)�Tf�g`e��2��V��)d�^.mb%��8#��Bg�b��vb����Q�+���K\���I'�P�W�&.
f�c������&��BR���o^CQ��P5P1|Ti =�I��M�L��_��z��J��ڕ�e����������Փ�3Z9��4Eݴ��e�)�i@+�)�A�8��0-Fq�kySf8#�4��F�+�d�ji�H���}-��TP��_3?dɺ4�K��@�C �4#J���4-�,#(Z�@71����Rm#N��$N�a����f�h_{�샛3�g�x�g�8��)vN�ҍ����ݑ�#���0M��f�BW��[�-�������e�p�����U/�4BZ:LQ&@j���E�H�����饻��~	�bi�1Z�Li���3�n��k�Q�e��}Tj5�RdU!b��)��r
��|�c�h9GK�e�B�����V@�0\>7�P!�ۖ���-J�~f����D��r��ǟx�
���LǢM�;���D���}�����<��3^�$��!3��6�-Pr����@�@���ۧ���@���^1� m
����3\��X+��jI��cs2Bu�ƺ��]�Jo��)[����{���^�k��/|���Mz�o�ar����԰���Zgm�v��M=�\��딽Щ.�����4]�FaD;��8�g�$���m��aڮ3�,�0H��Dl��$�-�J�41�!��f�f��_�I�e	t�4�?Kz��-Ys��bi�%Q:
#���mh�Y��ֳm{�95�63��g�<�O��	�8�>��So�r���hW6�wG�o�<���6�[KԭCo�Qc��h_[�h��r2���öh�h§"9Lh)��8I��1��0�x� �Ew��	�Ch���oh.Ac�+K���ں�R�&-@��8�S�[(��� Z"��\e�I&0V
�P8��p����hE�!\�w��2�D���E�nR�pH#��v�=ɭ�7��;�C=$�D[�FSb���\�88ë�>LI���&{�o=&/g�����v�I�1��,�Xڏ���.�s���x�"��~ZB�2-Xӕ*F���^DP�Z�u�?Z�1y�?�`���V�4j�+ח���﹥�~�2���9�a���0F9մJ�F�0+q�41�$���0�v���f�â+N���j��A���5�4c�jpM=��$i�[�$��
�W�T���J�:]s�*��j���Bx���c��~�z��c��M�������a���lS&�0ф�����:���%\\d�V���`� -�8a!��A�եUy�m�q��l&Xl�h��J��2K�|���5�%�Ҙð,)Y��.qw�R�S�K�#+�sS�|�"�ltw���X�b�x�Y
I��{	��x�*� �bS���
�)5��\+��la�Z�'��l,]������籼�,b(f��Alv{x��"�$yI6�����a��@N$��~ڼz�. @+%l���������ࣧ0�n��kK"��p�:t����d���lw�k���`�<�d�x���V�ew�]3C��������9��7uM��8���=�݂����)*~�d��i&�J�RT*U����b1��Fl��V2cY���z}�}�K_��N���l��~y���It�.�:��Ͳ�dG� �8����ז�G�>�kEڂ��P4��h=߀���\ݔ^!��4	3 �y엪�hY:�ǅ8�̰��-h�գ���XfO�+�Ӽ(J$��V/�R(�E���H���*sFK�U0:6Ɣ��쓣�� /q����RH%@��@3J���4�^.����f�|_fp�.�.�����ƍ��m��)j33��4��X��T�*��fV�f��� ���b���a�t��"D�6�:?���XYjK���-,�B&O�е;EI���,9g�'@�Cڌ&/3Y�[� ���O���_�bz�$}�=,w:�{�o��bMo��h٣%0�=H�8���R�\l�f��MM�@�z��v_"�(*#��Қ @�"���℺'�RE��T|K�]�h�Ē���`���D*�g��)fˁ�V*I@K��fot[=-�c��e���s%6��*�)�J�[&�b��2qL�� m4H(�ExX]�!�=gN? ��^c������}��El}DV�a��If��"�-��4<�O��V�\2�>ɜ�m��$�h��y|���x����;.�h�bv��O��6�VBw(�඾61��������]� U�k[Ç���:�gݘ/�qv�m�XF��l8�ޫ-�h�ی��c�`l���hY:v�yH���X:�x�`�A�L�V��r�
���b��t��z�tS��]����Q���(��2�!.&����1Z�y���Wey�X��B9���C��=�d�������Mc	-F�u7�(�"�
]i�c�R��s":#���E?��X/��)�̓�����r�Y|N�ej������8_�܂T]��y�h�JC����G��G��?~�yl�\��c=��@��_�L��T�@M�C������$�箶�Ƀ'+0Y�Ձ�Pgk�7��g	����%��FEX^[F���0��2H��o���-�����cm6�D �*�����3Tv ��ǌ�K �&�0/z�:�'�`�����+&OT��8���{��f��U�G���R�\�&&�ں&@ۨThikH@����21N.�R�dY)x�G8/y���8FЅ2����S@��u�qy��[m\�xӵ
F�6�E�q����sjz��YtG>�:�=��b�"	&$�B�r]�c�?�Y|n��������(�o�I�.��r�u���su���{���3֟��o���s��릾�Td��d��g~�)|�����=�R+[V\Fu�H�7/4�+�4
��������?����E���M,߃'u��Xm�w�o��Q�iIm�3�VA��Xǫ7��ǗVpy�/��LےiO1� HP-˘�Wn�e�Tϔ߳�\��$$�6��ZM͌B�@3@'��^@&K����m�ЪѪ|��A�N1y|�PZ�.Ru��K0�˨���,v�i31N��<[��^�r|G�P�<��` %�j�.`�	��K�aw$������D�RBws��
$�c
�_��"B�ǹ���]v��ͭf!�����u�̜KHf�����5E}<��PUo�ֿ��}�q���G�f�-�ؤ�(M���� P^��0n�-�����:Ѓ.~��E�l�����7ֱ�����hf^DTjE����1�/�|��O�i�������qw���C�� �=t2&���\��t�x�9�υ)�5n�g�-�q$b�a�׋���^^�K�4�װ��bA"�b����%	P�;@˕$�VjuGyA$�Ap%����H��%R,P�dY�ճ4�̰"ݷ����PThEp$�ӷ�4M`�7��}�-K鹽&c%��0*�z�� M}�)ӭ~03��'�ī,I�IG+���V�G��j0ϙ�+��$�t=^8���؂���ũX���(�v���>�V���{vA���׽���5�	΋ߗ���BM��g����:/ � fԃ�wQ��_�����l펃W�.����:.�RV�.Y��o�L,����>���?��M��L����N��d~8+��<�5tm������@+ۭ��q�uSJ�7:!���U\mź/Z�o�@�x=�ao\���b���1 �ZZTh��+L���j�v/�J9��z�M=�[g��x�6�a�XU�w���;�d�yL��)��2!�����{	�墽=_L�c�wfn[ݞ\�Ԧ�aX�^���X�H��b�V��N�#�Q�R,��d�2Cj���ߐ�0Dx&J݄��\MË�.3�ZY�1�}s��{�y�ÖY,?/�`Ϣ"y���n��}�� %�A݊���J%�+-q�z��\��Fb�P�O��l覆��b��f��_|��������Oiڛo��p�t �2a�?�e�<�d�_�����ݡ��7�B�b�@�H��r$���h=�p���/,�����P�,#	hㄦ%��._}s����2ձ2f�	�ei58Q ��u�H*�ݽK���K��9�ܰb;2��._�ۖ���XU�nfcy�I,'�ڦ�R�(�=�*��:J�*F�'�N,���<�z#�z��~���z�碽��Ë��&�$!Z�˘jԥg[m��QlLC+֥�LE9�F��ʬ�̹���>��Z�vwa�����#��9����{/לm��nAAK|�5�b*��?�3fg����(7�ڵ\Yٔu�KU�"�2���J�p��ŧ=�G�N�_>�iJ���M��=vB'o��\����}����N���@�;6QP�:H���}|��u����r��Z2ڵ+�=Za8c=Z�	",��t�-����K��R����R�{hsƷ�u+��3�)���:�rt�R*�uF(��,$�%�j���]�z����Yyݗ �%�e��l�q��a)s�V��K6��g�lԠ����=����Ëh-/a~� ^�r�G�����\�i]	��R;�|w��V@;n�x�>-��J��AN�ϛ�bޡtLA]�;0�j��階/�������C���ce����� 5E�!�6P�54C�v���'O���/M���ܿ&G5Y��bn�����������:��h�ӫ�J�D��)\i9ң}eisW阌�@�tA�
h�\�����ұ�����>���v�vh�h鱬����1���Q��V-��G�V��o���V,�a
4�x��"ߓ���7Z�f��ţ�#�O%N����իrq��H�,_��f���D'�8*0�5	��w��N���`vf
��vGO����1Z.DG�L��U@K!����;1ZHȆ����<����YN�@6��T��*߹XT�C���1�n!�\X�e�G͎�3�����_�t�����H	=�,۱�_,0]2�HG�����?����/v��ANV�^����@�����Q��a�$�ҶN�؇��� ����R��%���/m���J�%@�x~����--�v�G;r}���X�d�����b&ژ��xے���ߙ�s������f�v��Q�K3�ъ.j%�����]L7���jH��Z�g���s��E�ߞ9sF���C�m��	��>uJ~F�E�42�����0?U����x������񓢴�tK����םk����������Av/��	pkW���{e�u	�؇�hÈ��%=@�P�}|�c�p��^A��D:��@��1L�s�
6EM8΁���}��?>t��ҤG{ob�C�����k]�D���7'�� I���P>1`m٘�~ '�����-m��Ɂ� ,(L�m��`e�x׃@ۘ���C�� c,�AR�?f�B�ʹH������]����q����"�~�6?��@+Nƶ��Kɚ	<7�_�Vkł�Z���f��%������,QL�!P\ɀ�}=	*�    IDAT�Y�Ν;')Jv�_�������@���Cg���/a0r0}p��Cp����,І)��j}c���Nb��� 6� ��؟��"���Yqُъǵ7��Q�\��_��O���}����b�õ�1���Ǫ�����ӏ������Mlr|���W`���v��Kw����(�xOi�:�6<n�vMJ��^ڒұfW3���x5����KW�uP=*�k�ړ���>����Z���xZ0��s�4�HXfC����i���فZ�|�Ufh�{M���3�`��93��q�lI�[��NF*o�v7n�{��� 6���8<:>�!ʦ!��vc�3D�`´�:�̍�3�q|F����_\\ā�9���D�>�(�"0�"x��r�����M�5�x��9���F.��:+p4nZP��W������(���c�;�`���=���lv�|��fD��:ǽ�>�p��<����˯^�jh\t~��亳w>U�PO���J��x��=Ӽ0a���N69��
��+�����so����C,s��qyE7�6�$����
о��%�72M� ��Dm��HR7�ݐ^�8��Z��g�xj��.�2�m"��0̻ZI���� Z�1s�e�8Zκ�Hc�[.��˙{�;�|��;rt��c�)"$�¾3�`sC��Q�����*���AIp��nI�8��<�̳�v<{N��b	^ئ��^|%SÙ��p��%�6�p��9����6\X�~%�OF����#o�w�wh���H�"��}����=�0N�<��-��IFÐ�\_�KL�M�ҡ�X��:1���7�ɡMV�~Y��s�?r��p����"R~LY����-8q�Ȫ�>w��K�=��.�-s��uc�(�
��s��qp�ׅ̔`�-���Pf&1��=��Z�θ3����-U�{m�G��~�9���Z���<�e~v��fQx�ȏ���������(�����u�+eP�ۋ5h�zD�.�NR��#U���66%�o�є�r=G���b�A��ph� ���p��2��}��\�@kdb ��V#���;F����=��������0Zy��	]TL%8(h>>�������װ���(H<{eT�M,,���-hp��E����\�-� �����ݹ��=����gNOwuUO�:�ǂ�3޿_ę �2[]mf_�k��� C��n��'���p����w��7��Ec �Rr�Q]�c��+;���fb�w���ʪ �o{G�����|�W�����bo�sf�2�]ɴY
24g|2���"��P�iQD�>��eC��K�W�]}Y!+nw03K .�o8N��
���|
h�T��1D�r4����uը��h�
�+����y��Lm�B�,Аᒣ��N7�j�m5XAw����i�0�W��6E<��u؅���$�iTW�b�&�3��K@/��Q�X�{pb�:��~0�0ӑ�$!<�*�	��jK�Q	�1�͵�㹖A�h�pZN��H�G���q��� M��4���-H�wJ�Z��t�B�9_��L����`#0��!��������sؔ��Ka�0��@�>�V�*`.��l-���@��� �*T�VV�`�1Aw���+y����M8�e�M��9�X���9�C�c��Km��& #r�F؄�#g�&�h5�v{U�"w�(�O���i�f̰�A�I�Z#�SH<m8V��u+�����'GdwS�K-��!�u�뵦+�`�n�؂uՆ	mM��jT�ĉ?D������Q�+�4�u�W�Kpb�`��SA�=�?.v3P#n�c���B����~�����bc'��@ל-ҩ>#<�¤�?���#���WkÃ
N����H�>�E�Ń�2dX�&�dh�©P�禟�`v�f�=[^�����x!|*GU�P\�7�n�5�AϻȤ�������o��q�{S�L��L�*�BT�$S��?8kQL;�-���'�s��ݍB&(8�^�ŕ��pf�c;���w�XM�X<��!%L4!�sC5ǁ��%�IUD6R�JE��'׎$ȼ90i�#W�5f��z�6�
q�ٔ��!�d�7]��J���^�}�$��U���m�c@U�����ի���s&�jܝ�ȏ�-lA�I78O ���B��\8Js��G#�CE�w1��X���e��Oo��a#����]��@M-���sU^��=C�pk���E@�>���Q�~���b�v����w��P!�Er�ہ���&"��bc*&8a+\��B	�����?M��� y]L-,&;�m�B�yҢL����]D-�E���"@�yr�33���$��T=ԓ8i=�@��v����o��Q,�T$����$B���~Q����T�9��F�C�as��.�B^'�	�:\�l�%���5�nݠ�q?;��w6S�edg���옢�z�W���R������(���E$�[��@'ou��_���y��(��!)(������a#�2w8;�BE]�~3��~��m:���"���~���_�g��t�q�yҮI��-��KG�)%��ןO�	�T�d� �\^�nƲ*^�P�0F��g�m�鬢e�����"tU�OH��.��J����.;u�v,U�%���M���_�����p����܄M#�L��1��4��|��@$�<):6���s����~� _�� �4�)4
־�cĭ#>�� z�*����~�l)z&�Ħxc������>[^��[FM+��H{�d=/|�l)��R~o��A)��-���>Uo�\qK��#S�q�%	D��ީ9��!T��?q3U�ƶ�j)�Cq�r,�-�$�%l�h��=�~�JiV���k%������q�g˗�G����$�i*�S+���|�al1hN�L_�t�T>��1�Ӥ�rs��}�[���6�}���
=�6vtX�O�8�b���s������r��S�.,�&��eH6K�9<�"����#������!�֕/d�`#RṞQ�����V���N8F�
Â����f��&����/�_�.`�v�d,P�e&ph����Xo�&-�����s����t�x��hp�����Gս����3I9�Yɩ#o��f8I��x��������� ���"�\X ).Y"%m+�q�$����S���Kx�����r`UYF紘��2�;e��w
$�Gw����	N������.2��4�3mJ�\G����D����5�k8HK"mh�K�`�~��4�y�����T� �Ep���_��?�NQC�{.���c�S��}{Ha�p�t���.Vf9(k�8�s�$PK�fQ��NɌ�R��$Q�ȊW��T�O�A��#�#Ar�<cäC��Ҳ
�����Jݯ�L�zMB�����ֻ-!9����Z���j�fXI��e�ת��|�,�k�t����׮C�7�Uf�J{)�n�A�����,V�"s�G�BZ>,�ѿ��W�)�G:GB�1�`��m�nɚ|QUj=k��lN���A����y��ֵ�_��j5 �ko��\�=m�4F9=͞?&���M	ɤ���T ܅�;�q%`�9u"�.�r{�;p��c�PE�0hK����A�,1����^(�0��p�]<rv������A�����u�]*
A)���F�5ey��:]��T	j��m}Z�R��I�aO�iO<�K�2�	�	���!325GA����Y@'d�?t�8�����s"�����c��泖�̘뫆?8We ����\�M(�����boǓ$����W���I&�ɦ8
�����Ƿ���91Dhԟ�o~�E���q�9��I5���h����>���Pb�0�Ѽ+_ŭ�5�!���pc=�h~h)����/��i�篇X|߳J��L��E\k⇬�m�_��ޞڏ^���v�np�|���%�D����"!��Նwy8t_N	rC{K��&� �M�X�����*����2�%0�nz P�H�~�\�[>+�ĮɢYȡS�>d4���@fSP	.��2���y~O����/ �L��t�A���:��M�~�G	l��ɐC� �P���R�z�x��C��	l��s��1�u����r�b��#�	�"����'�v��X�P!���I#J��UY[a�ݬ��ܛȞ_�Q�o�lGd�KاFX��>�a��b�^�F�9����'>�0_U�B=�����p�',�d8v��5��N�@�b|���XU{��*����oW*�n�:۾
$~�<���d���	r�s�R���(���P��۞�g250�$Ǌ�!sU��6���+� (��sC��0�.��̆���g����d���a(��Q��h4OFKD��c£4��a"b�b��o9�`�O��8�.����P�Й�?�ŧu���� S�:��E�="�~f��A �gww�&P��NT�'�w���brr@tY�Y�%���Ҳũ�N�?HllXyX�v�uu��J#�ㇵ���d��8E�a�Ӭ�tB�Vv�E�����3�Л~�/6?�Z9�?<k��f�uI���Vxr�f-\��pZ����[#-�r[� i��K�TRbD��c�5�E���ߢ�\k_�r�6����� m�����9���Њ3����_4�A:\��	%?��������i�+[���5@�}Z��y�ម�
��g�����H,7@�g�e�U�LF��UA�V&ߢw�i���=z` {(o2�Ӷ�A��N�G�_>c��z�����hS��RݖE��A���K�����:j�2�C>b:���1uJce|cP0lqG��q�|QS���{GX�;�Ș)�\K���V�n����LJ%}4q �g��<ץ {Y��t�`��:mC�.��K��ypD%�Pm0�q�ϑ�W ��{��
�i^'s�?iqo��uo��V͓ңi�J	?������Y�� лi0�P� �r +"�#�K	�����J�Rআ�g�]U�2OZH"hE>,�(��z_ӔX"p���d�37aǡ@͠�ø �\�*ژSF��=�of�[K�y��{f�w���C�6��]/�E�3�cG��W�%�����̨��7 �3��#Hxw6ǩ����� ���E��I��I�P�gȁ���5����71���-�<���)u�r���iYd�6o�k�fslV�[��RkԓJ�
5���6����|&���A� 語��(�5N�mdd��Ro"I��5W��U� �D�,�F�p0��4�4*�N�vs���׀C��7��8���m��Q��'�	���\�R?y�q�;qȇ�ˏdmC���8�c�.fE�!C�J�1�a��dn�v�!*+�������hi�o<Ӂ�7� 2-��E�aFk�*�H��C<����K�
�����Zh6\%WaıVlTɒ=d�&�]�z��Hj�Ƣ j	=�b�t�����qlA�Z�����!N�:aoo���m��^��`N@�[9]H�����������y&�0TY���`�쎐�WU�e�j�%h��r?� �<���Η����\�I�N� ��k�Wo��z�ܢ�~��*�2�r�rr�������MFY�a�i\�|m;;x�.��%�����#��ӯ��)ۢc�-�(���wqA!͒ń)�T�9�f�1�t��U�O�̱��?�0J�P�S�*%=_��_��C)*?���~���
��|@���n!)����x.�tu)��`�r˝�V�L8�v��/dW�h!��''�J��\�vr�SNc ����� G��Z<eB6 ˌ�,�C{?ӭ�Xgzg�ֱ'G�(�BǮ2{,ӈI�����Db�q�(,�S�]ʲK��g:X�d�zhU�x�)VM�+��* �9Bp|�^i���9i<�����յ{��6�=�\������-�&�\�绦���b
*ڡP�瘚n	;��ش�*����']
�<��X[T+\j���`���dBc��d�U��/��s_�:�?�5�7�n�ot8�M��9� ��� ÔS-��&�ܤ�Yk�@N`�����qi��Q�"X���/N�DD�Dd�}��S
�����ms��"@..��l]�+���4>Ќ�I�g�r_M�B��0�&tl�a*��;ťL�"fYpe5G���)����{Vq�U��`GlSvf�	n��mP�R��Q�-�~�t9s�lg�X���̭���b�ךݫ�X�Fwͷ� )k��yg�,[��U�ު�_62�~��D�X#�6�ȗ�q?^}q��*��g�s���4��I����Y�E
�g��g ���?������q�A�
��U�|�/�R_ƭo9 7m4���[t�ˇ�Α�K(���:,)=/�GRu�QB�W�Q�T
4F!��/Na��ɬcD��̏i�V����G�P�^�5�ي��_&6����58WF��ZJ����S��;eI���U��~u0�UTkor�*5�م/�������#*C*m�!u�h��&��4��ZM鰣�&n����F�մ���O1߾��&yｔ�-�߇�SK�����!�d�w�O`�ʚs|��_`�X���cOr,eJ�bє0�0����}%����g��O'�s|�aK��I]�K�n�d��6��
�?�	G����"-ƞ"W�cBE�B�{,$�Ժxp�i�U��T���[t_>�����UE��2�Z��T��kD��c �����[Jd�a�B�i�:u[�������q7�pА�����	<-g-%���o�G�ԁ��7у���^��̰b��f�ě��R���x1�I��nF8/�h����q�8�m8 ��oЦ��aJ"���>�9˝��'�#RQ�ǜo��ǹQ;�y����&y���Tx|�}�h$(�:���m��|�K���0�폏J�U-�n�L���e�\�[B_�.�ꅑ��1��%[󁝛{B�"1] *�HP�d� ��AlmmI� >�
5�<����Xo���'��V:�tp �������hes���zNc
K�$	"1�S�6S���9�KnM�1�Zb&�g�I�U�ɻ=w�5v]_CaX�țT%���8Cv2�����E~��N��(Dw�cT���:!�,Ⱥ�a0%��3?3��vdr~Ҝ���/�R~��9 A?�$�Z7��J⚀$���Gf��S/۳�US�)"'=w�'xN�%Zt.�.�Ⳟ�"��
~�ۿ[���������͗�=o�=�-��*�;Z=M�����S�Ea��@-�N�x?9a�Z��
��ɓOK���)j��d���$�A��@ō"�� ��D�����p�a�9&V~�4}Z"Nw^�D ���7n��2؂�w�SNa��D����ɐ&�W}}|��8���Y]��L�4C����M"�s�q+3�:^xh��a�o?��h`s_tc��`+��5k�?ɽ>/��:�s8_�؝�N��L�}/�ēm���A��i'G�E�%�����k��ř���M���}ol:7�=�=T�@�97��Җ��=�}ꠠ_�uk�Y�M�~�.ۢ�k��&�%��²�WT9�_�)s�i	I��%ؤ����
��D?���8(�G� �z����uq<G�Z�_�z�h\��p����fH�D�Oz釺�#
�aD���'��dBa�{����B���6�r:�*K���[6^���E�
��ήT�Olݢ��+=na�tHW wI*�.���x�5�J_��a+&�=ۚ������_��@������N�ٰ�$;&�b�lsЄ��|��*�}��(�fk��]��� ��u�<�ef�:������ʝ��`4��9���(�q��q����#��c�O �a9��I�(F��"`��L$(i�R*"�'В��l�)[f=��܎��9�Z̞�o�Q
H��fQ6u8Y�fϝ,����6,�Uk~L�K����_���@P��rI�?��䝶�I7+$�?n=�r2s��<�ߩ�\*Z|S:\�k�k=i�G\H
*���R|��Z$7	lA�9��l������U��<��٪�8I�WʟI������
����� ZKy��@s$���);�]�1ve
�����ԅ������0�7��tIb؍q����
^�����_�(.�е��U��q�=�ݠ��Jg�$�?Z��rv�+˧�I��g�Frs��W�i�,����=���Ŝ�ݬ�Z��Cd>p��]�}*�(ggP�;R"�	/X�=����W(1�bL��i�Fr������,{��#j��2��]��3�n4|A�#�R���=�ܐ���vZ4K?b�6-˦LP�'���/VG-��v�=�n���5�Wn�b���H~X�GJ�Q^�X"F���~7�������z���x��B>]����^mX9(�S���G��>۬�iwE9aMu�L��[̒��X�'�m�%�ڵ+@���1��<���e����~�b˃�Q�5��T���+��I�oX/�x������:ޡ��B1�ʑ݋;��t���O	Rf��r�uq�d�yI�N������K�p�WF�D�k���=$�;�Vj_���ɗvY���P$���o��s��;�Ǩ�){����Rx!|�kG6�a�i�~Lc���P��_a9�Ryt������ɅP�:x��%����i�:m�]�u��ߝ�}�4 Tk��n������:�O0l����.�"6u&�o�����ؒ��t}��5S7>�9Ksq���S�r�h.DF(D"*��`�G2j^8�L�H�~��������2��V@)�1iAݿ������9O�ɯ�^�[���9ޯ{� ��amg+�ĮKg���B���M�E�w�U���W��ܶ��F�GJ˅.�r�A�����
��~~tB��B�٤���X����g�x[��9��?��� ɉ����D��Z����F�L�����)���,�?׏��o"=��2y�v���Js> m��A?���>��0jD}
�h�P��)�9�@Q[e5+�[��#�B("Fk�__<�w�Xd��}��0�@zf��-+��f�Pu��!("��B�&֊l��90��~m�V�s�_�	}zl�9 8��Z�p�0�co�j��Ԇi��%�4V��	���a�,nybU��=���.0�>�e�V�Jy�(K����{�{����PAvz�	D|S�[��o7hT��w��ɹ��Z�+$�"��:���@�=k���{k���ɴP0�a1ևL�;�!��;�4,�N6 �_?0M����WL� dS�f�dA`ɫ�_�Μ���n1bnT`د,�x��۝���sA�O���'h����Oa9��� ��7�Q��t��(���C0�KCd�]�?`�����E���"�]�S��z�SUk�-�)(06<�8>2�޹	@���=���7��.C�
�2v����50a5�'��{��(bѡ�	m̬kk/���J��-������4lbM���fP���a�E�����k�0'+٣���� �E7�-K���t3
je-�
1 �
qR?����}� ���i�aql��^;(!�w��#�_�x�Ԡ_�X����a��&4N�3(4�_ӄ�5�ĔHhU�G�ȹ�<��w0*6e
�"E֊���d�/\����`L��!������I��<�OՃ�4J�$>6�<KЙ8���U`��.Xmj݌�O5!0_�M��[�oK�3Ҳ�f�D�t��bԘC "�]k��Í	�gOm~��/�Uz�qk��-��ДPs�Ci���(5X`�ْQ	��u$?/��@}ל�]�����A:J�ߓ��7U�Ձ0�-MA�O2�Pا��:��CXA�aل����K�{�h�E1���%ڄ#A�.(��:@��t!�*7���[~ڊ�����X���礈��6�b��.�qkHܕ��r\]P���͟`�3J���V�%�[(����Np1�6��77hiUZ\F��A�L�L�ț���e���0�%��8�;��������E���2T^�8���W#Wi��I뮢Ae���`\��������t ǲ�ʴ�P9���Ѽc��IΧQtQ��3�l�%�~�ل�%�#Ǔ<�Y��r�˖�"A��I���Ȯ����ϫ�k��g�Z@�������ڽ�S /r>��?&x �먮��v���!��E�������|}���b��S�Є��s����U�?��L���fV�Ǚ�DN���L#Ylڣ�@ӱoC�����"=(e���޺k����ܤ����nl�0);#����o�W�ʐ{�hF��iҽVͭv�DWo������7.�J���-��]J��|8{/&��1����~����;v��ӫqHF�<N��囈������ĉ�V`j�8f���}��"4�t�>�	XAK����Q*��y��Z���+��A�J���\���~�XY�f����VM��\�/Z�2_w%��ݛq�����08ئ-�63�Z΋z�����jiC������POc��8)���L�s��A�^��Mg�k��{!�/��S��.��(��v�r��g��W�=Kh��Ν٢���J�����G�?�*�sڎ&�_H��eI�m���v�,��b'��=%��	�X��!9�q�8R��SI� ��S9
����EHSx2fP���..��#��43�K�g�dH��̧�ګ��h|����#�d{�)z�V�6�4f��b~�"0�Zwp�/5��J��@-B����	�۴w 4)�������T� X�=�4�J1�&�&ͯDb�F�����7eV�v�����B���F��b�1|T^� A�H-m9����Kn��)쩉��2�]��?4~��wMe�*�O���|�0}X6��e(�P�>��poϹ��˛ [���G�� i��iJ�O_SJT��;��/��b��4�MɌ�V��=�?J�'�<��Rz������	�m�r�-��?�s��� ��>�v��Qo9/J��:gk�翘��n�)�1uÐ�*�킚anbS;K�[��f����=\Z��΢4n���pV�F����	jQ����Y\/��>�:c�5��1�j����/�\|fNKA��de��ř��+U)�9���'��zi�m�O9P�9������4{?���f��S��HUO�Uo�� �Hu�O��l+�0O�gpv�� �MS��=$��4	%y&�"|�A�_C�CF$���B@�ZՅ�Wǭ[9��m�V��P+8�3"->�9`AY��r���
�';W��,5�s��a��-<��z`�����l�	�,�̲{�	��D�#����Z�~��(_��^�9��-���|�S�ԇȎlt�w|�����q���0�rD~�=������b� 8��
:�h'�����+�Y|�M����Il�F��
�>�1�����,H.��t%����r����=������{�=kd���q�ՑVEi�(3����L0�rP�bz�<�a�,�b��ֿ@Mɟ���^���EY႘�ޱ{I��MW;��c� ZY�����-D��mɃy��MN�H���ڨ��1�����,���$7���z�ռN.�dxZ�qG���?�����I!8թI�����}�ʞ%͸AD�K9�%7n!b�g��6}����G.�M��H��f%�k�+��o`�����*J�eM�|P�
ӵ�I!��m�P��J����"��묱et�8�vpf�91��ɩQ�"Qe6�ҿUx��9�=�6�5��;g�wp�S�M᭒~�{y�����=�ɵ���vy�7'\�b^��3V�%��T11�^�w{�#l����}p���`��ø�/�-�����{�35�>29��0��<2��ИYۄj��;/����,�[�������������8{��A(CB�׿\+2?�%���S�;&��˫t�Yp`mʢt����n��X��$D�W�' Eœ���=x_!Z�JoP���B"N��s�9!�kb���<���ISD����L鈻���Wg�a�$��R-+}��W��q#1�9?|T�8�c��ķ��fO%{�d��:��g�7�n�+X�����u~3��T?��^�*a��N�᷾�1���xq��b>���~���ֻy���l��"+'ׂ�� <�^'Q@%}&�t�Ƣ9좤Y��7�� �GY�<�(<%`G��qK4��Ύ�֟BA$ݖ$Q�]Æ�`+�L��8j)�9�h[��=Y����SB�U�+5�غћ��D���o�Es= }xm�Á���ɠ��HMDK�c�o×�3�1�\�J�`R������p"xAO����xlXŢ8�jx��g�|�d[��L�{���Ï�B�C)���n�?]���^E+i�XX�����c���V��������7.Z
#Р(���vv&����v^È��RT*���@�j���>���+���3�z�s�\��H5��[g�0�s�T�N� ����u
������:s}O�*��p���,o(���,��A�VF���tkij��$�;�/�J��s��/�h o��I�GE���8�kM
]���4��h��9�h)������Y��xh�nH��KS��|t�Ky��Gk���+��XV/�Oc�8m[5�����4z>��?�aE�Y �g���������	�͉�Ï)Ü�˯m��p��{'�Z�\'�Y���73 ���efh�p/�<:Ȉ��-;2���E��}8� �h�w}G%�xO��X��@1����m��7�=5H�L�M����}s#��w�#��G�!��C�p��́
��`�����A�cD����i�s�io�T������Z�9�&�(~�5���\��>�ND�RP�&�y���<�.V�W�-{���/��L<�����b4�)\�h��a�Ȩ�7
�l>0��ȚD���#���%j�'�������l��͔����P�R�kZC:���˿Fc�2A�Gbo�Xg�������e1�M�n���r%�ba���X|sQ��H���R�!������g;6��ĳ�܂S��<t	��qI�鞅�!C�i��Q������ 49P�e���NXo~ݝ�g�=����0J�p�&�fTt���2����>]��_�Ɠ6k���ֹ�6��C+?�C���i�<"�ja��A��R4�,!�e,�E���γAV$�J��1&����P-NP�A�v���!����:�]��9^��ݻ���&�+�G�:���S\e���f���Kk-I����-�\ꎛ�����*�g^��&P<�)��dJ��O |�?ل���LfY���x{��(�����k����V�y��b��o�F׶��mL\��߆� f�c���Sfs��yԯH�Y��4�FĢ~���r/��#L��8���98|�@Pm������XT��3�؅�K�FJ.�?d���NK�����FhGr�*Q�nθMW�񧨆'������}�u;��?��p㯎=M?htMÓ{�m��Q[��it���i5>�Hs>�): �H�<p��V��ܒB��n��u�6�"#��h*����j�`syo{7�D_%:�6Md�jl畗p�:f:[�-׸�]CQ�~���[��Q�%���w\ec{<<�G���K���$=�s���.�n�ǩK:���7�rE��D��� �
?/��O�{��Ikv�hp,�a�1���Q3)*�$�Ժ����s��ړ:" �}-U b6{�7;����+�E��n��<3�ۺ�FQ��0&���F8-W<0	�<��X��Q�o��4�2e"8�n"��z��'~�_��Jk��C��g���]J��/�)7�}U��2�v�
� �C����掗5���hi������4�w��x^\�d^��l�=ր����G�̕>�[�Xg���~���"�A�m�^����M��.F��2P�,�M����*�������Aj5��=�y*��0T+�j%����>�T���TnOy�r���G	pLc�P���@�����@���nŚP�c�.�I�t������`�.�\�"C�*��� ެ���ܘ�̺����:�$B�J&�`�L���ȰP\��?(���W�0P�1kVEC��s$�f֢I�=�󸛆�y�����m�K\S��v��Һ%�7^$�8����o,A��ԕ��=K��.��?�,�w������w�Y��)�N���PAMc��V����?}ڟ�6pK�^�]�Hb�y>��ѩ���0]�o=W�,2c�o���}�����]�p	�h�}��p���mW���9w��\�yj�[>�ъ�,v���7#��������ɹ���:`�N��g��;H����|7��MD�B���\�5F��1���R|���j�A�
E�ٲ��/�Tr↌a��bx�|�Qi��N������.���޸�ot���_��[�G�׍����̜a�EV�Y���6�b9��-a��~�t�_�b�:��%��K:��0 ��;�i�z��k�-�Z��
"���Y�oV��2�7�=$@�����YV���cͶ?'�S<��L���_N�ϡ�������٠�BLt4苺���-z�Y���Q��-0qU�"�I?�� ���Ǌx��M?�8�Q`�6���3kD�$A�4��{�}b�@S����e�9|�r-� �`tRQ\ke�Q�!��bs���p_�p�`��J$6�^��n)���bT�H��
T��M����.D;2�����]���?��Q��]��[�"9c�W����Oa�vܼ��?L�v��:����Y}���%����6���?oR\�Ògc8������s
Z�\y��4�v��I�Z�Y�T*�|ٯ�7Q���A�w�g��a�������������n��*O˶r��f�h��݌��qf6~1�zö?\���o�CP޹����qB�c�h8����I3�S���tVSidԀ�Í}�V�!AE�N?��j�+���ݻ�p�]��,dM�����w�ZL����"�`}Dl����XZJb�ad������C9{zcEo__�s���.�X��Dʌ9��m8�W�Ƅ$�����+Ɍ���mx��bUx��<�e�5NĜ��.u��a��[�)��Ђ��T�l'��`��'�7x}��]�X��~,�K���ݨv��i<��������l�Jk}��ɷZ�yh�&@x���D����+E��"&B�U����c��݀{Q]v���e>�;�_�C�S�\N-�4Oc��w�g+�S��N�c'}��d��{X4����an|��L�Q"~K�C��s�ְ� ~�q5AM�JH�:T{�����D�ZUe�P]����ߩ�9������;|X�=�.X&������>���>�H�5�M��6{J����D����N6�9��u.��G�lM��d.Z��λ:���l����o]ťGsb�F���[`�rȄ6��v���������r����,'}E����g���G����*j��0����R����N�a�tÛcțs�1�"�G��}�6 ���r�&.{E�񴪅š��?}�O�o��R4����R��{���~�w�[��pS�vw�s�ސ�9؋���x�;�W�r������M�Y_d2�d�?9m`d���]Sl��C��"��cʁ�(O<��8��D���.߷�*����Y��FP#���!c^=�HYG<eY��5YޚDl-�X9����X���d#��gK
��Ī�H�$\�=�2�*/��U`y�B#���G�?[՗*K�2����ݓ�e�e[��l�UyKd,͆�،<ìa4M�m�7V
�">$ ��TV�H{kd�>�q�dD�]m��-Z�k'>�:��E<y����x�7,�	�'�@/�g#����S�����(�8��N����ϟ���<�H��]�J��")H���Ď9p'����������!�ؑ�D牅ܫF00C��"F�A~��غx��(ӄ��>*��M2Aౚ�bXZ�69_SǔV��P|�8�z\�H,�î�p���R?)��ěG5����7?��U�
�
��	�(n/d��5���S�!V�S��ǡ�c>c�1lb���^yTz����Zo7'���`,��6.��]p�]��H���߬?2B(�SU9Re��z�*�(�@i�FUi\�ĄsSh/=��կOqo]O����bfH׃���m\���i��r}m�7���Ջ43̘`��%��H
���'bٟWy��(��cp��ˊa��J��? �m!6sD=��d�D�����Gc�upʾY��d����Ϗo2,<�t4'��X��sy������/r�Ź�?�W<�eٳO���`�JY
/��3z�TS�%׸ƥ��-��w�<1Y�%�$z�3GP#��<�"{r%��ŋ!�΢ �.$)�76lB<�"�I"������O͐�W������O⪨#�F�`{g3|�#�aQ�-��Q��F?�[�p޹�>Rn����0_���?J���s�2mU��z�ؾ�뺝33S���%oK�b�|NsM�5A��Dxu�w���F�_�WUt�ά��uQG�/B���3�ճ��a� *5&�+վ��v�R����{�	`E�Ɠwz�ˇa2zy��b�F�l%Ĭb�4=XJ�U���M0BRT�X1���vA�,d�����ƌQ	V�d��M%V�QNrő���H Pi9��g�
f$F�c�o�H}ؐ���7(��5<?�F��/w��R���-��N��}+�h3�y��=Ԙ��7��H㼕��ޜ�M^�R��;��*���ou�&�^�p7��� Ї��=��"xIpSN{|f���^���$����V���Yk����>e��,���/��dJy���� ��툑�(o6k���d��5�YyQ�,pS(�9+~��u�W�Ȍ��e��P̤ia5�	Z�*� 3�U���F	�Ā�d���j:�/Pt�6`�o��2�����t�ƳA�HC	����ѮqwGh�I�
>��P��d�.I#�����6���ZW�{���rr[f>@f��6��-{X�>rI|a-�?��++���W���n���ԘQ&x~	�9W
α����ˇzp�͍i�r>��S�tDO]d�wnzD0i�7x�4���{�!J^�d�O��#C�'�T��Ɍ ȣ,��G�[�@�b3{c��ed���Ki�\Z�S��-nt%>ةUjl����4¯����y�F}4a��E����S-aʱ���>GuKI�:�eT������RJ�����B�8�q�$�@�ׅ$���3�I�L����z�t��d�Zx�[	������*�G6^�D%�8sѾ
be��[�frk��֘��8A53k�� ڧg~BX�t~� 鸯�����i�eg'Zh���kBnD�����������{ۦK�A:����@@B�F�.�f i�:���a ��~������g���������S]��V۹�ʱhr<N�j�gU�[ӻA�:F"�Fr"��z�B���Hz�+Q.���x��GS�h�ZA��H�_:=|��lȈ�㓱H�(&fr����i�#��S!X Zk���&  ���MA!�΄("G��("č�o�ǧ6��K��l�����ߢ��,� U(�U�W�Mt{�W��nY9�}�j�G�a�h��)W�Dc.\��3�z�ۜ����^($��N�DKxL;GɳH�%���3�c|�_�_���W��UX��� T��"�ق��X0�h=��,l`&��O
�����}���8~݄��{<����-�8�c�|M��{���V=�?j�~��}�������c��� :�v��M�B�z\�Y>�!���/SN�_������Y�Կ�F��4�r0I����@J"-($�5�ĄEZMp��� �x�{x�_�W�a{�2���2h�"?�:ȿ/,-���(Y�������%�c����r��w��F�Ȕ!h�s"�å���8T�(������ G��z
����b����n��2�xO�]�"��]�ps�5���*ۂ�����@G���9ظ$�el�
�h���3B���)�\���=y"��ܽ�b[�AȵHQ�����S^W�SlRc	���K�α��uߐ]C#�Ys�v��j�@)�Z$*E�)~�\��MP�i�rn�;*`{o ���
~��A&8e�m��(Pg �O��\��z�;i����gW�)��J55�,���Dʞ�5kG��F�Se?d"�lŞ.�ϝ��(�r��]�m�~����-�4IH�?H�!����Nh{�\��2t�����$2~��?�M7F�醽KƵe��6��NA��Z�G�#r�>�R! W	��
��x���pZ�7^��a&?Zj��"a�~��Vuԟ��Iޮ�5��-��� �n�}�=x�`3D:2���Ys�|�pE�Ki7�E�<��v�:'��0�_��,���9:Bc�m U!!�\S��2��y�I\�VLm�qH��K��Q߂�Tټ�E�g!�
����Ҳhc�(Nӱ��0�^�{J�L.CԿ��b�gĈ��`�m��'�E��F����0L}XM9U8�;٢I#����ehS�N�����&��E��C�|�%(�*g�َo �z�>k^� �_�{��:���� Ϋs�8;2.!94�#*:�c1
Q����y �s����ۤGI�P�~Pz9K���q3l�!��G�m�p��*��[����J�_n���x0��L�b<�4l���9}0ĻMt��1
��?&�l�E�!U+�!8|c ��ӂl�*~�,Ǭ-�l�X"�)�T$儒�>���\4�|e��.�5m��S�&'5���o�\Ŷ����д�G�&�����Tm\�׿�[F�f�QWZ����@�t���m�f�xCv'��P���u����o?)I-"&�ae��ǯ׵8�yZv��va�M���� :!�s�2ݵh5��Wl}�S$�7���	��O����|�,7O���R��������dO��x߿�B*04e���K����ɧ���O��qC��c���q_�, O�E�����π�����X�.�{��?���T�'���k0Ğ�z��Jq�3̮y9C���t�3 uD?�i�a��}���]�^�5���`Qz������bT����!��=�r2VA�ۂ�ق�y+9=~�X�O���#&d�Q��f8�o��&S:r�Y(�8X�Y�R^�v��O

jZ�1�'��v���)X�\0��\r��{ɋ�h*���'^xˡj�/ʠO!'o.�@]w�?aA�Ev)�K�ϗ�y4m S�{o��������ߍ~�řQ��%ە�WB��Q�G$���}KX�N Ʒk�ӕ�4�&���e�2��PG{-�X[L�t+�x�A���n��6�R�a�ȘAx��;b�
���v�����o@ ���~�v����iǀt㇝���
yڄ*���Em�R6(��6��	O�=����� ����x�-�X�����J�^��ާ%5�ꕜ�H|ժ��t�\k�����Ր�Rj�A�!���"	�%�mP학�Nw,]��N7R���T��ht�_�Ot�e���P$�]i��aX����bi�q5"s��D��k�����Q�
��c��ѐ��3�y��#X |�l7��*:���f�23`DŴ��g���Ə>,K���%~h�3�EJ����B�!�U�e⡊CD}����E��5c�T�������,��f���6�q�% R�h֥(.v���V�p�D��U�(����I��
��=�v�嶇"?�s8ʱ�_�Aj�5`	(.,ŖLD7��8�>ͯoagQT�TNw�3�AZ~s��|�m:�����J穤T�W/�K���$p����#>��^�uNp��@#�J_d�R��8T88x�jA��IE����s�[z0�d��J��S|�Ulp�Mb(:�)��9QIs!����g�V�f���9J���Ҿ��2l6����n�&��1��nJ�u��&%�M� ���������@�A�!�~�Qyf��w���#m]_��(Dv>̈&��f]huhM>���m�'\��[�\~���qL�*T�{����T����['��|���C�'S���aV՝��gHs��>��f��+�h�QZ�w�+�
~$f.S<��Єd�!�z�
��L������ ��a�������D�ƥk^�Fh���v*��o�͈Z%�`'-h99������A�8�#o�`�6ޟ��I�
�&��2�O���N�$��)t&��e琓Ox�tyl,���,�¦N�� l눙�Ƃ���X��pj�:&q�
������u��L��8�2����{��i� 1���x�u�T�0�+������m5|�S�I��S�1ƎLs�C4�m�j���8�S�N��j��d�%	D�@�Wc3�F��}\(���,�zI1�LD�>�0�j�V�.kZ�G�����~��	�eq]��<������&O���b��,p{j��k��%��c�����C��CX��/=��xp��(-�����!mN�!��˱��1�;�eulFF�����;�L��W��O�(:%�{�-&(ڵ����dtF�l}�V�#���^V�ǟT���N�!�\�<����Llb�t�L��F=�w�j�7$#r�A5�&z3�b��"ڵ��֋���릀������Ǯt��\%��kGɩ�G ��C��%w[�P#��~`�lO�V���JGK�Ԛ���Fz��r��&l�xV�]�{MZ�T��{;���d��P���[UV�HMi�J��*:�=@c�P�Dfz0k�(��2�
h���;D��w�>��uz��{�zA������K_�/	�\x(1���嗓������R;'������v^dzo�$Ӏ芺�������u����2��Uz���x5|	쩘�A�S1�5��:��f_d��qZ�@|��y�}�w��H�{4��[^sG�\����٣�y��@��J=]�m&t�=2U����qh�t�fH�t�,:C
("M��`�����'>�A���i?���J�����-E��~e��xh�vp�%~#D��(��H9��$SP�z�6��bˀ�8gHs�ϒ�	r��~�a�%��db���ɟ�����J�v�G�I:"�
���y��/�s=և9Vс��-y2�,��z�Y�z����o���;��o^�^y���w��T��@8z����F�\�~��E$�.O_�?�a�1!��c�%5��[�{/�o쁃i:,���>��/ċsu�m�e�2��i�{�����#˽�c�sKud5��u7%�Ȕt9���=i�俕K����8�� IC�l�U�D/'��3��������
�>Q5�_�9RW��]�{!���F�G������]�6o'���M���{{��i?	�@dVp�`Wi�=�nF����_a��#Adm��7FL�?^͉�%�w	�˖�9��bX%��e��e�B�U<�f��v�Zx�����а�2�]z=s'��Χ��~�I�C�&tIv�-�N:��9�S�Y�?�j�U?>�Y��v���5�l\��K�W���N#�H�=I1�@�vM��L>�������2m�*f�č�i>����`���Cz��%
�Do.�j�D?��>J�����ΟS��QP�aF�2�3@{��g��d$��jU�-N/��9�0AzLI6c��f6��]z���Fl��&�1�4�}���)���n8��$&.j��rr���Lp'+N�������G����z�������pd�|e�t��K�&�I����憗��}�D�����T�&Q��!ǔ����Q�0�٢?s�b�UC�nI�F/�)����5:`����4���ݓZݠ�hؾ�2�E�o�ł�/y�8
�q��m�N���*7��$Ma��>��k���{�Ĥ�X�x���.�\�%����T����d��2+,��,��᎔̘��<�@O�27�%��TѼ��em'5н�X}��4� �/���%)xE9)�Aa.��ۛTb�&0���Z��������@������Q(��ܟG�=џ	�x� [��-���M(+n)��Z��ϰ8�t��f*�R'2a֏��2{^"�O9����܊5S@����mV��hI�$({9kH̑�@Yd�U���v`k��!E�f�<��+��*�|�<�j�(�#��{��b��B�W��ـZ�YUNy�/^���Ԃ�M�N���g�`@��]M�U}P���B�2��3�Ԛ�8��O������V�L�wX���Jom���.0��M�We{�O����-*�gnl�2�}N�,�u�"��י7֣�)Y+�(�|��7$V$��g	�C�xr��d\����P��4 Js]�MmMK�e�c�)\~ժ�H=g(֘ՠ~ :Ӈ�n�?��2X��L.bVp.�1�ch�))�i��lp�h����l�$��ﲥSܻ��ڑ�V��E�����9�ʽ���$##B�K�Ҳ�ܢ|���,GQ����ʽN�{2(��e�e�l��^⧧\��C�77,�i���榩%��X������8 UD��F=Y�%D�1��8��Y��7�Dyco�Ix��-������H�6%����� J�H#���ۊ2��>62��r�����Tק��A\4��VR珣�pl�����̞Ip�����/ۥ���&D����QL�/xw��d+����"��Y�IG>����1z�����&q&�p�����y�|�1��
w?^�i��V���<�n��;�<�w���A40m�g��GNf�憢�F���+c��Ä���S�Z���;G<��8����0�w���'�yy S����p8������K����ܷ�*� �s���t��OH���CG�'� "���Pr���؞3F2H`�ۻg��`���m���X��u�Yh;��O)����G�環O�������r�] ���,��G�U]j&�1-M^� }ws��K��X�R��4�c/�9B��v%f�j���`��(��2�mX��j]�ö�+*TVљ4ʩ@�,�@�]ٞl|-�nRS�0�9M҃5���nw�I@ڰ0���j�ͺ��2����r �>b]�4<������h��259��;ݤ7y���U���̧6.^lϰ3|3>�7��|o<��������NН\
�a����\e+z�Z����@�}��j����O
o�������v� ���İ����ň��Ò�Y��A�V�����z0	*�c���Dú'�sԛYH<ɏGFqѦ���$�T�M���.�-Q�d�Z` d�A�����^&oe_^�e��yL�Kټ����������)G:h���o~��}�衪�LMKK,���a��]K^�����_Xm������Dǀ7o��w�%zs�_:��xĊ
]������'��%�)�=�:%]����.�O$��)mv��Q&��],@�KyJFM7�d[���N�C ���)eV�pi�<#v�>g\h+�!R�eո��л=�oY7�:Y�=�R�9���������|gth�:��&��W��~��O����;�eq�l�����E�?<l)j��i��~�O��t��z)��L}���l��[Qa��gۯq�0�/�w�Q'
���(�p]<����M�E��U��أ�um6�t�6�/�f$h��8*XE�IȌS="f�&* �LUh8�p�fP�-�Y��`�?8H}D�	���D�"�b��y��@rh���h6>�d�=Wݡ�h�{��"�@��*,Q��Q1���t�
T<��������a��V�̰i��gz~�w��`%�!:1^��4B��rmH�������C��da���ȝ�ͅ��V�ܲ<���3�k�:)�2�\���_{��8�R� �� f�d3�=�C1Lc4�����w�d)f+�H��ߟ��;r�"E�{�G�U;ų+z��)8���ڞ?��8����	ѣeJ"ي�u��#=�(��T<��{<Z-ԝ
�4BHq���W6���z�b��#0ؗ�S���������L���n�X�+�B��J�6т��������ꎱ���$6�Xe�<{���v���Hy���ɫ��C+��$�ج��	ئ��W�t��~�U������g��'��4��~]\�6q�W���f���WY)�z{�^w7���<p���[�	e���_���� %Aݳ�L%��v�g/ш6u��J�X���m�G!�Cy��c�xR&�T
vM��BtH�I-��s��U�f�a/Ep�=��da(�`y�i "�a�	� +�VLv4`Ĉ����t*J�q��>�T�+7����h���O�g��D�\<��O��`17X�d�\hG��@���Ȁ���%+�ɳ�@�\���v���^����#:%�{�]�6D�+i}ǲz��-6}���N;>���vڪM�Θ`����FK���1�؎<�'����t��h���i�z��I�8��w�N��}z�ш�&;�@8�k����"i�-��\m\>���;Ps��e;��WZp�:��穷�0��v|[���A/lBE��	B��=�(���(��RϤ=%7�	�<��.�U�<�o��ݴ��%�b�:8�0X��X6�G�4b��ׇ�4Yr�Te:�ӀD�Ƚ�W�JU�������^9՜+uc�1h�+y-�&/d��=���0N���EEE���%&&�7��uiz��a�������1�T���%+RDnL�5�p(�{����L��KUJ�D�gA�]�Si�
 �EY��T����YB:	�vO�uj;ʒJ&nYu%t���E�?�$��ww�ǒ�ԫc5$ ?�r�O���V}5P�mv�����8m�3���<'����w��(�>s�%��E\�ȩ3�"��J��E��"�Q�Z�K�g��+�7��[%X�1�@@)�)��XP,mL(UtjU� [� 
\���争�Hg���F��_��լNy����'<�
��)cYg�RS�DZ*Q�y��y@��3D���ʗ&�PF ��8��QQV	j�bG��𜸫�4Iq'��B~JB�]n��sC���?7S���<��=���7�х�����t]>O����l�e�[�m�K��uw�Z�����>v)=��
�mi�,D�q�k�ׯ"���l�&JbaXC-]sy�F O}4�!�|)W��f�6U��"�[���1�f;�n������'��)y���EYgN�I{?�ե��8z�F�13+w��������I��vҞ!�#s���9���,�Ӭ<�����DN6k����k���g/�y���_����9Ik�0`��4 ]Rه�C�I���i܆�����`�3��4�`Fs��.����1?(o*@���N5���x!!Iϴ�A,d`f�) d"Z{��~�|ȏ,�0-�1ӌ�zi#T�!�i%n�8h���pƑVð?h�:�R�qp����&��v==�O:�A��#y�y���9h�l�V���x@�e�M)�9�-�wj������ud�G��
о�#��UK�N�
H��8���W�Tp������P��������������� t'e�f��~�?�g�@^|_k5v��l�%��Vt�Q@\h��B4�t5,�s�4��ETQk^��3��k�#`g�{2�`4����R�C�gxi�ju�*�TE>ҭr�u�aIʖF\M&�0$��M�9@���T��_����Q4P}Ы���.��|�]�����t7'i9@�u䑀V=�Ө<(����w��0��o��G{�q��n�JWPH0�J��LR��%`Qr@ 	���*;w�SR}�^�oR3q����G����.��#PfE��xd�C�v#���/��%�yNH���S���|��
�tӂ���yUw`{#E���Ng����Dv&��9���_����&��a��Tt��"Q�v�u��+D��;^`�<d�O u$�mu�U�v�vS��������+'�㰡<�p���W���W��4����C��-q�	�Q��H����)�����Ko͝8�I8��2�m�V�i.n��4t�`����<1��E�)��~߳����_�)8Q��HkQ�I����Y���߆|�`��v)�m1������0lGPѨ$81��y���_� ���c���!7������d��X�7GQsŶ�l�[Sd'ȫG�W���"�P���rqh y���3���e�oK�2��c�LYJ)n9�C����$:��i�~���6��1H
��wPd�Yxb��f�(bh���:�l�Ě��E���7�Q'\��w"��G�Qc��m�a�U���ː��g8��1����,�2�d�DbH�No;-������8�H݂�jO�f�u���6�з��6&
��i���ٕ'33�;.?}�z�]"(CviA����kI������R�(�#�?�Ʒe=����l�_�!v���GwT�$^7�<�4I2W�4�NM)�	�(��|xv�0��6<�ʈ9�^�obR��:���>����|��|o��H���(c^�"\�0@�,ک���2C{��i�*��������_[[B&���! �`F!~w�a:^JI�4��e��L��~���@i�G��9��!E������Q�2[o`�e��PzO��΅H��{��y���w}�>�����u�~>Vgg�T.SiwD�O�Mm���T��\�SQ�iY��4V��92��b��1s?2P%t�#�R=�r�d��h=[ F�%ӑ�fFg*�ySn3�Z�q��7Yi�Ep�Vv]�0a%2�^�n ���.�e��P�}�߸�}��!ax6�.��[:���)�f	R���CC�FQ�7`l�z}�[8��U����<`�]�>L�=a��匽���$�QQ�ZL�U���c�qS� �Y�d�ܤ=�F�Yҙ/M�.L�Ʌ8"y�H���O(��ոÍ�ۡ�]W�)����#4@�t����]�N��"�j�F�!��M��*����p����3��3����֘�-D��EN�������:/�G�g�aϭ�a������	v����[���y���4�M�B�C��ȥ���cR�w�qʳ��\&2a���V㓥c��9�CQD�S��Z�'#-$m�kr���
T���	ʙ��*q�����$�B��V��\�B�����r��^.�[�>��)�97l�I���==���6,{m�0�Ⱦ�$vT�<X+���55��i֎�R�u>\�2�]>7�����m��2��Q���S��59���ʽa���Hd�O��L��TNJv���v�I[
i8��E����l�1����ݔ��f=m�8@z��-Kz<e�.��� ���K�ک�Z��?�g�����h�R�����9��9?(������Z������O���
h�Y�>6L(�bI{�!�HQ�!�A�}`x5��x��!���<��۟�}����x���^U����$m<G,ʔ�������cm�h��A��>v��Ѣw�(��Al^�P�p��P����Y$�{�v76o�n�p�Ӫ}s�v1l-�q��Ǒ"��e�Rg�lC	���v�g��)2D1vͿ�����/� �զ��ի���
n>�?0ؽT#��[���Vt�1E���w����0��anӌ����]��<�?W���GJFHcM.�R�)l���o���#�0��o������[��m#+��.;�XE�XB) �G>��f9%��h֖�e�����-�y{66�'��6@I�F�
��<���PZ��P9�Q���%�g��z=ǧ�S�p�qy����O!�o#�/[��|�yK��=�U��/�y[��'��~��j�R��/Ī4�0����ܻ%������!U��c4?�J�a��>5���4������kd�|�&�5*�7v��t�y��E������E��
p,�ž�����(�w�ԇ�|���ޡ3��9��H\i�NUs�ad���!����펒^����h�o�8{�)	���.yE
>���m�)�į�U/(�l�k%���Wz�Jw��eG�j�1���C���@�� &u-�`�x`cV�Đ�6�R��5X�Y?/��vK��Ө���;yO�(��z��71�����g����z�;)��Tq$|����Y��T�.L��s#�S����4�����_TCK��@m�hv��I^�c�?��f������f3� ����6o�|�k�I"?=��a�_:k�{�� L8`,�����U�'g��;����-ˠИD�ż$d]��
X/M�VD�P���%�?,��L���GGn��-�����_��q�}T���r�ӭ(L�{�w	�ǋ�6�J����'G�k�R}��Zۻûl2��ڔi�t�B���Qp�K�"h1$ƭ���p�o��00��ƀ��"��c9x<��~A�]�bi���S�f���s.KW���6{��}%1$͓��k#��x�]��P9-$Sz�!:��մ0Ul'�]��2zí��N����!]�Iҟ|���nrJ-F�yt�4����~��~�7���T j��AU��.��R���.цnZR��Fs��	�)z���j�П�w	�I<���u���0�������/�{�j$��5���*�%���1��8��\㿦�-aKt{�j�iX�����pf���)'e�~�c S:�3#�ָb�Q�⒝���.\���?V�(z7qaz�c�w�b`L'��P�%#,����n��np�^���A��ʹ�����m3A�-ڑ��.iMCKd� KC�܄Yׂ7ۈ�T]����2E��_���i/r�Z�q!ٷ�s�6����_�",��,V ߍH�6��V����S��>�5�]�1_~:����uc�"Ud$3��r���
Eۼ���o�PV#L�����2:i֪�{�q��Bʦ^�u�_T��s~W�ys�"��᠟�ܢ&͠�=~[&m�Wd���v�?�:h۞�D%���ht$�@wd�7���+QE�n�k�7Hq��Ѯ�s���r[s	^�0�fĬK6+��9g3��S'ck}
��Y4ؿ맀�� Q�E�G�ff�f�2�N�z2�O[��5��چ�#��K��=��}SoM�zd�<�2���GB��2P\�Ҽ�i�-K��7uWm�9R�G|4%�l��z���p�/}9���0���(���D(��$X�wS$�@s/M��#�5\'�,�(zM��c�g\�;�@���ǽ��E.�Z�OZ���R�D�����i����\�S�:��p u�~��S�B�X�B��HP q�����
�݆ ���D�z5<u��C��%=�I�_���W�8H �.�͊i��;�ӯ�E���/$�R�!8	f�W%�	Rq[����)�����-��^��Y�z�$zje�/S2ӿ�p	w��yc4�(��7�cN��Ҏҕ
}��5��xT "�Xl�X<�����{X!�i��z�;}����cA�~��LS�%f
��u�I�u���'���� ���x����o��Ѧ���&X�
_�f�M�z>��Vy%>��V����<�I�m�$��τ"'`��޹2
Ą.������N�{�7.�8���&.�D�0:���^�c�u�S�-���Q=r➔De���pE������fm� qς?(�"��OO�B��X��V74|��{�)���1�9�Y��Ό�e��1�����-x���_D"�NYuVs�f��ﰊ�?>��ր:*ƧMO�-� ���1�=z��R2��5=_YCQ���ؠ�I](��.�E��s�i������ꓷ�Q�ҕP�[�5�4}�	w��T�ۿ~���.�q���Ѿ&�C�~��O��Уq�� ��`r�?�W���|��#�~�8�NT������ow:w���⹁�^�������	J�S-X�kv�J���@�����hl��3���Cᦣ��lcMl����GT���o"�]�u���U��A�>��Z$hXk��j��f���G�t�)�7	ِ(`	�g�S������Y-��O��l��'�7��>��q��xT�@�V��M��=�"7ۋ��6
�渾�����7P���}��c�!���l-����i���?����u��~��$C�]��R;E���:~Pd��C��Re��oQ�T���S߮�s��Ck�)�P0�4�0���� +"0.]Ӓ��q�kv$�X����GU�&���~ߐf!rёB��O@ꐈ���]���m�O�G�&"�z�`�M�+M(�[*��R���Nxp}�^�U�z{ڜ���8��tc���������䘂�.��*;�6;�)u�O�~�c}���dzW���"%_h�eI�\&�a P��=�3i2�5��Ȗ��h���zK�tE.���+)�"@�.*��,��t��Uk��2�L�����w���9#�$<���R��E9L՞O��ן��5XSm������i�ڢ��0/�ݳ,�/,٪�Z(L	�`?bm��ڸ��h���W�?������� A�Hv2K'����+c������D�/^����'�*�B���I�a�������Z2p��Ϩ�B�9߼�<�^i�,�8���_��"��=��co_^c�=��$&2o0�����1-Bp�.�.��5R��f�iS�@봗Q�ڳ�O2"X��CE�c�f��B�:W8�;Ǒ�>��w��{AI��[y�ՀZ����B���>Q�� L4|҂�m�M���[�dTd:����@����CNT���+o��k$�I�o�̡X��FyIv��+�,_:ﻔ���r�ϧ�Y�<& �n}���Ҥ�Z7y��E\e�gPYQb�ɇ�_Qg�L�ŀr�|{�,ʎ���f�|"{��цW;-�:y��L$�Le-�z�P���a-fTbP�,�E�#T���Bb��ׄ��św`2�/��h�d��G`��	53�%����I���\�b�_��4�-��P~�������0+ueF���B�I����yZ���;���MK/�qt�>d^�y@���w�Orf�mq�u���&���0HpZ�&{�>���t��Xm�'[��b���fg�xx�����X�F�U/�ng��ֆ��� A�ᆓ=)ȝh#d�]� k��`���R~�zV�����a��\e�o������OR�8V��
|�۠暠����� �"xO+2��k`l�F���9�L\ߒ{՜߂�Nudؠk�U_T�#��T�69%��+F��޻��)��n6Fi[	�钧��'��~@4ļ��d����d�,��QJ��M��c�R ��cg/_�L��p�Υ�w#��Ji̩�bb8U"E�]�?7��Pm����r��0��C�ܚyg@�o��q8kY%c�[A�hlk�?%	t%042� ��*�t�˄B�D6*HBy�Wற���GM6p}����8����F��uOom8f�]	r-qtwf����9��E��.;OVY�y���R��G����bR�5����܆�R�8H*n�mjH��Y�}�]�d�E��� �g� �*�>54��ܳ���I��b�R6;�4�	8�5_��������CT߸V!�E���r!���K���)M��󧭡sz����$�tF,�|�~3���7���q�ʼ)6��G~�����7L�@|a��*ˁ@��蟭 @7=�1��.�_����N��-�0�6S�X�n�G�xS鮝OM-&�Kߟ��~t׌Ȭ��S�����Z�ޔ��n&9�0�75k��S�I}2�={(�=�J� l����dl�RYy��R_�H�J	dG��}�zb�4ҥf���D�xm�pS����������,-�	�l�I&�+��RG�l8HH~I�~���Wn��*��T�뒵�ם6V�f�{ �=u��a��.J��yys��Uϡ@1�(F+��!N���q�4�晃=���C؊��;�Ċ�_�bS]:p�ꑯQa�%#ԣf %%%�
�׋E1݋t��pA�ŜA�3"�*聟����e',�޻�a��(�lp�K�� -G�5T�&q���@$�y�ƙLj��F ݐ%�N��|�]R��R�]�����ʓ�fK�󦇠�L,ML	����j�Z�)]�]���F+p�ZRH�}�\�p�O����F�x�S�εq|u�� �(�Oa�	.�}���*أA6[��F�J�G��p��~|t�����/ws/���DgEp�g��ZV��jnG��S���4�fM�LA�ddj�Fϫ'�ݹ�`�8$'��w��<}��/"�FBR@�2�����菥J�k���!@=��K�tU�t���[����=�
�Hh��Q^"�(�$�'.���F��t>��B���r�8,�2�|��r~%�<�3�]�y!w��7��p-��ݯ�f(**k:b���5��DT��GFF�>n�2G))���Z&���ݻ�e�TH��
�	��mА�[��$o��X�	��i5��q�r��s�WF��*��*ۖ��ů���v��x?��|x��wV̰羄��_��q�{K}Ip��t������`��S�N��D�nOz�ԛS�@��VJ_����<��A+\P����?�Ai`=���;����p�w��(�R��o '��s�^�\^��j��)k2��Y	E��Xȶ̡�^)��i�{vC�G(�OG�TLib������
ċh��u(_m��W�T��������t.�O��u�n�	�\_|S��C8�l��s�&ijk�l��{0���
�S�Pd��-�8e�8t�����W�
����[�6��Q3[s�<���y��\U��P��D��s墅�1��CZ�]I������yp���#T1�*�tG"���L�^����B<���>�6"v��`�W2�@�G�|6�^����|�S�ȅ�YSl���LE�Hr'ʺz����?5= ��3x�|^:.���ۈ���\��-K���ƝTs5�A����H���
j��+�X�8�W[$�H�����v�,�F�'�wSB�Fy���V�71qs�Z�<�F�8W���Ί62�z�y�ܼ�?s;�s��|]m2��{�el�O��M4��*A���6��+5�N޻�w�J�"�U05�gSYe~^����U�A頿��M
�v��`D�nl��w{�E1_2�-���H?J�Ǘ��h�E�>j4�6��`��S������-������N�|�ͦ"p��l�qw攓�C��'��)�֯�Fv|*�ߖ���CXUIZ^?ߔ�'��8���w;mN�)󧰆�_��_�|6-�q��gOG���{G���Y�?�XC�i�i��d�8ݥ.��Y�yN��������I���*�Q�`g�y&�	�.��������2L��pߺ�`X�ʂ�j�&y�P�����$�-a�~Ꭸ�,B�$FT�8�)	�w}�{��e�Ei���\F"��wE�-t__*�5�����͖	�[ ���J`�l�MNC]����ҀB@��\ȗ�e��cJ���O�D>��h���lA�g`��#.tY�f>!�K�^ʕ9�p�-M���EK�Y\/q�+(�K*)Cw`T�ί6��|���%d��X��A/�a�S~M�U�m�^�5�#�-�EY�!5d;�y��޴>d#�ۖ��`u�E��rt���\�5}Pzx�Y��h�V]�Fy��x�<��?���+�&Z���e� �ݝ�������,8�tp'�38���;<���}��������gU��P�&P���p�;�!.~`�x�����%�:�$i����G�V^,�;<�پ��������?���Nt���T��M�c@��A2[��@��6�����>�+^��R-�LEs�O��3��59��( �u�򷶇��)�뼜k)���M?�Y
8O.���҃�����l؄N`����m'*��cM0C#Y;{��=8Ê2�K�^B>������'6飸��n��2�
D�,�YK��ɳ�I��ѦZCe����6�Ț�B.�v4��VF�:�W���ª����
|�	j��H���Tb��$�=�#��X`��h8�s�j���� �l��p��F�Ĭ�:�de8�؉��(b-�+{.�AC F_/�� �P�{�/_�F��1�{�T�חoN�eq�l?�1`fv�=��z����gm(��ޣ�M��zAL+u^�@��Zk�tǍ��E�,C�WK\E+c��J��o�ʝ����<$�Ę[���J�r�0A���1�B���pbA��<�*���w�����No�>����E(�}cӿ�K0�����.,]/�#%16�O�%�(�饽�h�2~a�/�9mt�)(��0c+������O�#�ļ՝�wn�kZ��@t�~+v	s�V���";�V�����Yi٪�,0?�A�xP%�ם��tUI�}�o����Ɨ?�暭2�s�
���b˘ə��A2��r#�A"��p�K}�,�E{�'T���g�zQ/&Shf�t�5�S6wq]�z���1�H�ɓ톸"@8%	pA35��Lɑ���t�!�PA��:J�lь��ߜ'䓶Av)���G���t$W8N�YǕ�ܛ��8����Yt+7f~_�m��^`�i*��hX����m9�fJ�B���f%G0�5�mxN��@7(П	DVUV��GV��s*����D���Ġ�'��ʏy�����=�Yu���
��C�j+C.D2d�;rI+`�XKt�e��?	����@��_]������n֞Ď�!�*6���
4��(���Q�[0j�P� �e�檩���BR�Pv��|��|�<����v4��J~�S�HǴ?�}�*����lG岨$��7F�fT!(�|*q���3����WD�'a��B�7����Fi�>��O3���u��]�M��������ѵ�\���y�	_�� ��3t)�柤J�{T����))�d<��-�NFQ]C9�S�o#k���5���n��?I�q�	CT��K���w>��#�(��X>(WC���̈́�h�?��I �G�EP�K	�%s� �rx�y{Kz�N:����o�)^�$���#��$-B����?bs�:Y���WE�4&��(_1|�j	0�c^���hm�zQ޸��#�&�#*���%7r�-��B���n��(Z���8H!�o��8��f�<-t(��<�dN4k�:�t�ې:��7��D�)�mKfO�������,ߧ�JfGkF�r)��s\�������"ޫm�RT���,��)�隔�ʡ3��8q���OZJ�JЖ��x�h"��g
}f��s�!�އD�=r�~�V�J�`�9�o�v~�l7������2�X8��x���7�y�Ųl��@O�	&����|S�=M�U�P�=�7�Z!�,�����:� �H�vIn�N�wëU �<y�<��0e8���!���aP�&����v�3���(�z|��O�ɷI%w|y
xS�?�R��u��vW2#-�B!�,��KZQuU%�f�<^��|4,݈&,}x!��2̧4�{���f��)-�g������Hw�>�p�w�;������T�����46B}�l,_9�7�J�O�&�B6���C�[w�<|�:��\���wó�S5��_���;ŕ�T?c2��k/��}�3��k`v����)������lj"�LEO����P�y9bf�ٴc��Z�M���|�o~�0�P������.������[wg�J��;�Z@#>���
�w����+i<�(�e�X^fD.D8�|:I��D��z3vK�3I*w�a)!�e��B[W���� $(Oa���z)�����>��4I��+����N��f��ta3��Me�y�Ѫ%��m*%���g���R������"51�gü���jh��~����ʫH]ۮ�~;�n��h���L���M���~�o4}ZM��}a%A�_�d>�%�e�mQK�?}R[��T�$My�G�_�����#*:t�}��k��e%��PLء�S�-�,������� ��T�<�C<���S���>����gT��E��f�w��k��
�շ�����Lj6t���"IagI˯0����S����g.t�j� X��="����qB�@H��FZ�Y��?��M�,��+����i5��Iz��� ��Fw<ig���دwP�KZ��i2���Z����d
�#B@}ֽbf�e	��s�Y���s�ϭ�$�:DB�@N+w���W�F�ߖt��!9B�ve��\�(����%�w>@��	�a�|��۽���2��_>�{OՍ�~z�-" �x�
�|�j�xe Y�,�ׅ������DB����	Ah��W��_���JmTN>��g	�� c	�?�S|8���@�"E�1��Wn��P&�n&t���i^-����!�7]T*ãSR������:���r�p��V���bU�:I��4Mh@�wVi���cv���Mn[� e��{���t�tsJ:�!J^c/��h�44s�W��!:����5.Q�Ѳ�O�ή�O���p�.����ٙ:%�����D���+c,8��f�tH��m
�u��r{��Z�Y(곭l$�4��v̖ ���U��q���o��Z/�� 삟E0,���~�Ie��B�����
4���^�Fyn�ܜ��>�OOy�Ө��`����g�3�-6�Uo��U Я�<9�yWY6��	�</\�z�  Uk�@�9���3htu�lmR��$�0�-�iY!T�}������6�|�@��!�򤒜�D�<ɑߒ�Qt=���o{b�;���-"�?�o�y��$�O���ϻ(�OS_N�>D�WX �1�pĢ��V�jV��p�˒_��D^�[������;���H�]Вl��<��핉��*Ǜ`�h�O|<?�>
نl��o�>��g�?�v�JY�CwMc�a��	ӭ�ν�b/�U%��׃����B%�3�p�෵_� � �m�ޞߎK�\r�9����5>i��d��L1�p:_݊��e�K*:�?~Ē�db��yo�{�3�,�䠟W��{�ŀ4��.��Y*�x�=�t�����zX>�-:�jW���M�+eˍf�}�/�%��>��ܰ&d�?�z�L�H?�}@���iEs�Ƹ�"�t2�������3����#7)[�|3�������qd�9��]����Pg��Rh\��cc择�7|�@�F-29i
񱁼Jy��x0	��j�fT��P
|�G7![o����I7d�n}��ǵoz���6���� ��eoGmjWK��%Z�\�)��1Z,��T��s;�ӊMA0�rX!�p�G�rR�'�����+x5��C;V3E��w�Y�2�4]!9F߿�������/`,jYT��=���"�x]f�%���'������D����uE����v�3������SK;ĕa7�BS�����T��1g/�ܣ���O�+�3�_p;i�#@e��Ն�,�b5�|�qɼ*��P���v�uME�UMۀ�u��4�'G���s'��슿M�ȵeɲ�����4�xP36�ǚ�^�8݄w��=V��d��F(I�XV�Ѯ&}e��7�!Z1��i�bJH#W��c��cë�c�"���/7"���nZ�L�;ɗ�x�n��qS�~�@��R��*��CEv�c�eE����5I3�V##c��	=I)�
6�%?�x��ێ#�,Y�Y�\+�~��Q{M/ cf��Sbd}�df;���c��̪���
Re�=����P�bʷ?�����Z�x��1��OqCQ�'8w��j�hn�BQ<6E��l���Fu��$�W���wХ׍*���d�G8H(͚�ߠ���4j\rq��_hd唝�Hn��sY��{X�U�H�>0���^�t��ݲ	�m�)*N���9l�ݨ��Ę(�\���y8�l�Y@�$G\GI����'�{��g f��1k�^���͡_��w<��C{O��ϥz䝯�����2�da��
d#S#:���gp��/�2*��Fz�x�>�\q�GH�k��<{����Zw=w�C��$$zxT�.>쥠��W�>�V��+���� n~�"8� K�*��}|��l	a�OV�W���c!�3C��7��9�S�m��=H��X3��y�'����.޵������>L`�t�d.����w��ϳ<�VB����2����ԥYw�#p#����'�8���z�� �T���j�q΍0��*RY�g�7���w��sz�e9=sNZ�C/OyᏪ��Fi	//�](��'7�[�F�	�	U_�	��8��8�p�ARU'����E�Y��-(�+S���q)�%h�>��bNP=�H�Y��tq@ �h10 ��<�~��9QiTS���]]qcV~u���0���r�t��I� ��7��J¤@��מ����G�2}1��Ĳ�%�;Oy!W�y���siQ7v(?I��Ҟ붞ש��h'6�J�H@�ɭ�L{��ۡ�+Ɵ�'>�e���'�Z��]B�L%�@e>�^#�0[H���e<�8��o3ŀYz;�[ؗ�+y2��r*��s>f�M_��#�oβ�$��e���e��?�HG��s� G$��4n�p�UO�ۻ��}�Θq �B��j��M�	�da��j��~WM^�H/�H���p��*Tc��0��~>��5i�[;�_��7{i�������`=��z�J�K���Bb�b��*���r��^5}�$4C��R��_���+���%e+f��Fbol?j���]��p]0q]?)@�/@�Ӛ�(&�:��⻝Z������K���Vo$�+[$�����atcv���N����v}����'sS��E��a�Mĕ	&����2�BJ��&{�� SxteEʰX�%fe2(�����aN����"�9q�iRny�) �����7�0�̃��J��7=<�7!��Ήا$�#^��q�7f��������OQ�7�qs6����,�1�&Z(W��+_�
gû;�X�)̂�K5 �s�Z+!����n���¿�i`�{7�p�B��j a�da���i)?�9�<t����ݕ8ȃ�!*Z�S�:ν;&��6k�LD����f��Ϳ�>[B��y��wI�Bx�'_���mȤ�g-�n��҂���pؔ��y����Es5�z��kJ�}&��� ����sǩ6�1��d���Cp�x���5U�[�Lj�Y��#��>D�$!Ayj�&v<z����$� ��1�4?mM^B|��c��'cJ >�-���GS��z]+N�s����������r�&/l}�.����,������,{\��&��dh�R�j�'�p!�L
�	�i^��a�`r�i�� ��&Y,�ޔ������Zgj�zd��ke�|c�ڕ�("�V2��鬘&i��N%�c���͏� �WdYWS�2P�c�G�9"m;������j���h<���#���*PΑ��zq:v" .��,t�܎ܴ�}5&_~$8'R���SI-n�~�ì�.��\Ք�s�L�N�ټ<�b�;�6�s�&Y�;�Ѡ�#9T�~9">z� �*���)Q�4�K�\�V�#�1���<�%ߌ&e�h�tUP��ﺏ�� ^�nW�ݐw\�L��eG�I����79�f��ᓏ��6& ~h<�dM�ɵqL�M�IE���<�"�A=@'�*X����� 8�)g4��s����qr˜	�.��M��? ��
��hb,��d�d����p�{�4;*���[�-&��M�r6���O�
�Nײ�Y�H*��%Mf������yS)��D
���t1$o$���dwu�=)Cg3����������{ �ݷ�3V��Lř�c����l�վ��I�kJ�n��.�'GFMf�&2�m�M�� ��������~��Q���(B[�s��c��|�-򎍉μ:�W��ȍ���Z[,������z`��	��w߯a ��ܾ�U�&	�=��S�&��鴘&�"��+��ˊ��q1>'��7�(?��A;��'
�� `,,���O)�H�kz�A8g"�l1$( �-�Q2�QG���� �"E�fv�F8�Y�J�,�@tW\!��,��i]9��ne{�Zz%�t�q��8��~������y6�݈��iț��рF��:��v��i_G���4���SؘZ�Ro:�b|�rV]K��`o��xj�`Q�-�F�~�V}��HeJ��FZ�J�e�)^�0P��C�R�/�&�$Pk�h�����h�6Կp�Ś�����fX~��CT�x[�vf��kY����͛��|�NX�We.�v�J��V�~{�)B HOam���X�	183�c��o��zRi�
�[������+:k��vn��tZ���2Ɗ�,�d��)��i�$c�.(�@M��(��\��# .i�����^|����;��)�+�5L=��w�IC�����a�"�j]*vZ�,V->C}�������K݃@��i���Z�_j׉o�3�o�܁��1�l����w:��R�OC�ϥK�H_�HH&�b���tvn0l�Z`�*:Q���N���� ��<	�xߟR����w��tO����������%��s�Q���z��iC�NHH��ә��q�,8V��>�-!{�'�:|Y��sX��%;"�A��R㟃ˀ|L��h�F��bL9p״i5.�U&M/�ln:]r�s^���,Uמ�n��9��3���j����[�>V��Ul��ӄ��:=��D�l��/���\�q����|=�������W�jz�`4e�U�n��2���؟���d�H�	�lJdK�%TH���* N���4}��ǹd
 2Q�����ڏ`b1���U{ZcϚ24�羀 ��}|w�ѱA���q�Q���\�A�qnNt�^�:^�f�g�`��b��?ؿÈ���T�}�|��P��PSL]6@e��.�J�@
h�9�1��OJ�:��a�ׄ������D��CIW�B7:��<�h�_z��-��^��KKv�2�}�~��u
>�������6��1iի-hXS��,��u���WZ��D?��}hgG-\wZ�@LB�^����[�<�P�0�#o>��f�o�`�g������E�
�wN��F7H��%��Ư$�V��it�:TZ:x�4&��ݺ��Hضp%�G�wf�U�S
�['&��>?���4�c��q�t����;99q���8_�ԧ|�Zw�a;@ /�3�ʀ���F�.��� ����E�������x�I�QÞr�?o��)�w��?��uCmxۙAID�nڡ��Ȃ\�+#(��������zV老-+�&Nt3f$F��\l�@e%P� W��މ=U���*!tJ 8���:�N)�>��@�ِ�] 8*ܵ8�)�ey��N������)�3)暭g��i>��|��1�&�8E���CԢ�iYc�Rj���G=p,#��/&�jW�`_8�ac�iu��%�g8:ɛic��{>�y����I�'҄���f�J��Z6��r���/�$z�z%8��-w��P%٥Y/˧3�l�(��%��ƫ"�����F� HJI�hG����E�^��wX���м������"*]�UG`$���O�u��m���K��}[~_��4���h#�s�W��>�J���ڃ�{��n.3z�|<#��vnn�.���^�����5,��Ifvw54B�,��2����G�����&DE�8�"�pP����L�� 4~La�ިB���7�K����s�n�o�a�i������ke�yi �\�E4)(��Q��*yK$������9{:���ʒԽ��9�k9�gxx�Ѓ��iJ���(�0��0�����$㭍H��c�@*Y�m�xęv}��`�� LUcXY��s/[�8s�J��`��I+�*��ko��,Z���a����O�z�Ā
i�B9p�ib�\<�Qaw�\�d\�l�ǎ�i{M��.��_q�v���`�l`�|ʉ��z�O��m�K�ْ��a�\�/���Ȉ��(�K����4<Z�؇��á�Ni�k;�b��Ð��N����W�J���G8���,W��:�.�@��[�>]x}�j=Ξ��C�C��
T��8|�E��Lw+!>y����Q�Niσ�z"yƉfa�7�tp>v�)aNY��o��{�t�;I��,c�vk�ԛ0�^Rg�<�ń�%ee�yqPu2h0��f��Hx��BAT�N
	Z����]�����jK�R�ۦ��r`ك�fi�2�#5^1!.��1���"'��\\M��	�hg�@�O�Mz���Z�ՂT����7�֖�h���+���2g�?�� �\f2R��?<�L2�&�	 X�7�S#S�FB�V�I��L<�Q���G�kw�m�ǽ��5�Đ\��������|A�@9�����,����3�rN_F~���ԧ����w=�z(�j�٫��翑��g�<a��A7����6F ��}���-�z^��*/OEh���ds>���D�/�3Dxi�c$K#`����	4�iV8�b_W�t��,���-�_���g�×�E��iϵ�]��9�1vZ�~ɶn�T�|�L�E��mD��֨
}p�ux'�D�e�$~e� �坜�x!w
�J�@Ϗr>���B�0�̐jF_����B�h���8 �b��BV?1�Ռ=^�����`���,�Ǽ�I� q���UL���&B��{o��'�
�����\�ҝ�(��PMղ;2��A&��FW�>l'��C%��;����ʆ�?|�`t�R4R:���b�Խ�y�y9WT!��'$�d�5�ũ���p���?�L�]�y
I�?��$��sF� �Uƙwɑ� ��KVԬ-�-�~��K��P�A�H����7���7/��_��+_�����_̰hյﱳ�) ��KJ
��ؠ<f�,���x����(!+]F�ڤ��ګ�K�M�K�Va�NJ�͝��R��I� W��@]��"��ͫ�^׏!e$gs!יM9�m�ov�\V�q�[\M�?����X,��j��G_�kCk��~���x�V8�_��"����r!���2���́��HϮ㥺����R��˴�u&{�]'�isL�$�w����YhJ^��I>6�)+nA�TE-�!a�^3�ے�8�r�m=C��
����<4��D���@�}c�{Cݘ`�!�l���V�BF�a����@��D��C~�om��o�5
��j�d<��O�.҄�ڹ�B�{��Z�$��{̔�_��s*Tr~�X���nПs'��ĵ��;]Y1������}�7�ql��nϵ][S�Rrb3�iB�g���1C��+���d�ǅ�<�9�β�b�2�9mg�q�UH�`�����J>���*Ԍa����=H�mb�p�|R�f�4�%Y�t:�YF�/2�A�p�ˢFJ*t�@~gF��$2øڰ�5 �9�Lyt� ���E���>A�ˏ�搃�"�#�A��<C���^��(?�|��Uk�ڮ���LmMk$Ge�{�:��i�,��H
"�:�-V����t�	�� �TK�e��G�M9�a�_se�7�q�����8�ʂ�-�`H"�i(���F&�B�gR͠o����β��0�%o2�'���@*�;�ʘ����-����I�������(9�
�H��^r���x�x�jv��3��y��_��=-�P����p.q~�w�aª�&��*������0�]��)]7�T
��P�2�n�a�Њ���Ә8z����L30�p$�� ϭZ��z){Ο��2RБ4��_es�{+@e��F˃T�P�-������5AL�+m�|ypn���)J��@�A�!�����q�}0a2$F�z��J��q ���yk�߶��ʾ��dE��Z��Q�v��w�@���`h�|D�A���d,ȗw��C+��wnE>Ų0&>���%�xw)�a��I�_��Ll�T�e/J+���ߠ܃��ꍩ�)����jD������lG���q��_�r>����?�,���]1��xg�p.脂^���: {/s��&?��:�of[���"�I��(m]�s�8?Jv��ޫ�=/�Q �����-k0&L�N���*��\�B�	o-PZ�ka��Z,��4�����b&҉*Q�͕����@�(c��_�U��D�w�mK�Ɋ�5�g��ϊu����?V���9�#Ц8�TЊ�R-O/�+ً}䪣�|��^��,N҇'�4,���k����f����A�\���?+n�@�u��7���F�����7w]/Ñ���\U��K��7���sh��a>�U��P������}a%̆��7oI��$�葆���![b���	u��VPb�4Y�N��-�y�?ճ\�hC��w��	�G�>E$ �>O^�Z5�fe��*Wo������lӔ�/~W�l.�*��*aϛ�?D�{���][}��f���c|��a��@iN���\�K{��R��w�foJ�=����d�C�?o-�1�"%��D#k ?&���P]n��i��sN�Ei�d�shL�?��S���y0�ׅ�#�N��q�����7<�&���>�����(��ky�!џKt�9{���8)�|��g�ܷZ��ǰ���hmD��@���4lP�T�}b\��}��)�R��c��[���,0�z�>[(�uI(+>��\0����i�ն�M�zA���!R)���{DTv���X�3�ˋ�W���j�o>t�s�ʓSk`�fl��B�ގ&�7W@y�IBn��gw<8y[��(�/N�n�L�}Y#�-������biY���h�i�t�N���TZ�v�z�"mF`\9m��%X����*��?v^����5�L�8�.7�x��#_�h��lBa�:���Ӱ(�� �b'�/�i�"�v������陻YɎ�}�Z*�zD�h�&���>���?��$s�����z��%�XA#J����l����=�ܧ=����N�����6f�SD��e��ќ���8��/�m���a��������^{1�F�󝩁��ú��	����U�.���T�[�h���VUS���o�_"�V7T�Ҕ=��¶T�2;X�9*��vb@'���#wpݏ��GA��"�j��_ͦ�͍�y�-���Z�Ļ���^��TD|�C�+A_����u��꾈�PW�QF���(��9ޮ��V�7����&��n�1_�aꂆ�,����[�A������5��]�����M���A��"�Љ	t�Q<��1s�.	�^��N��b���$
uMѧ�ڣ��;WD�zh�X��.F�⭇�e�Yri -Z�눿КP��_�C�"Q!�A]�O�61ve7i�`�E�\As�Ms�[`	,��	�G5���V�F���������h�Lo��A<H��r�A��Lu4]^t��R�͊)��稀]�k��k���)�,]������Q�v�����`��H��׊����T��D���oW���L�M]٥����u[f�B��%���UT�Xz�_Y�Gr��g"����C��R �[y�.�|F;�x"|��s%�z�!�>���������P�u5Ã_�=�����t7����J��~Q$�nf	Mp��=0~�?G^�i���}8I�s4�F~�?�q��S��EP�w��
��o������h��r��Һ����_e���#�|(��=��x������l��BS��DG˻#��t�?tY�"tN� 5�7ᙖVO��X��s�	�*k��Ɗ����������H��vf�)�I�nZrS���wC�&Չ��~���Rs��q|6c�����^�y�\^A����!�C08���2ܼ�3�.!>z�q�͎�;�>�^��h�3m��+\�F��L�ީ�ݞl���~E�!���f��U��s^�Cyx>v0x%/Ƨ;�l^��6T]��� ����v�:>��S�t���)9��K]�a������_l|�QP=KP�t�2����(�v	�}bdg�޷�X@�j���.!������A�柺l6I�a��9��m~���!�|�'4j��:YC��� y+�UJy�{z"=|?<�W��s�����3�ȦҢܬ���(�E���V�^\yD��R[��k9�fY�T�~���p8�����c�;��v�лu���R��]�;�H:���V���/��P��6��o��h)�J%&F&l]�|���<�Dn��V��ʠ��� V�� �)����Z���������Ɍ,�~g5l����T)��^y'V���L,8A��<'p�²���Y�OCL )�2�{�R=o�#�^t�Q���+-%���W��H���L�`F~�UM����X�)���t�M靟\�Ü�	+�x�Hm^u���q�bʚ����Et��/5QnCI>a�4h�`�*B,����4qDOK���VU��|=@\���m~�/u�u�v=y�2��>��I���<���:�y����Օr�=k�I��b��C��66�A�Н����$9�K�,y*a�RR(���Fi�߆t̜5bzR�_��9Q�[o�T��-o�����m���;$����˅ƍ��:��j�� n�=�"�7+#)�Rz���[,�s�qW���F��G�T2����.2w���D����c��r���)��X%�n���I�� ����%�whݴ	��FۘE��s<f7X�qH�����������p�ݸ� �&ڢ�Y�����i���Tҁqo��{��S�|ܸ��uLG�9 �������쓀g-ڦ/-KB�!V�b�ȃA-x�3�?Կ�?{�<�It���+���w�,�R��r5�ZEt��葁N����zƙ0޸Z%��
S��b��h*T�_�"�#�v��O�u��śQ�����ōL���¤-[�
��ñ�T�?Y)L4�q{Ȅe�/A��`���7�8�S�nR���Y��Z�痠�x�{vk��'W3�7�'ܷ��T�N{�i<K˔�n���B-�V���]ݕv�%��4e�$��;��L�3��H}W�|��c�h`�=>�M3��f�e
T�����$(�=�/����l���ǳ�7�.��n�|</qn�����WD	���ꚉ����b�8�	n����L&=/V�T�I)r��Y�kEj��˧K�: >B����%f��Ru��DCdF7*�r��b���H_^E˪�by�=�����,��^�K�`�o�>�ۿ&#��M~h���8-6J!	`��k�~}c%=T��Nۉ	����� �ĮBgV~%2Z�Ol�}�?�)	���][ �|�[�[�l��æ��ʹ�s�$�g��5�����lqP����<ִ+dV��_]�=�Q���7Tf�b��m�iBR;@M���'��菃f�#�k�W|���3�o�d�+XK���%�)ngj�S� )G��]y�B@�VĹJ�N�� ��(,M�_9��(|-
|g��m�V���݋$i�Z�����5�u��g�5�bB��R����aXo����l��]�7��d�(�U稷��B����U�y���b�����2q��3X[MG))/��m���g���U��o�ݜE�v:�:°C����)g"��Q'���c����rՓQ�{ؿh�x9�����x]+��p|Q����"8� S�J��鱓p||Y	�0�3yꉌ_]z(��P����/6�� ��g�lH�=D�� �����\BӋqS:��jQH9��Ȟ5��װ�V�ao�D�Z����#i�5�<x�w&�Z���aB+JS\Iz���wͭ$wܷwV�i~��P��Is��*""�c�l"��X�AZjH�`~���Avkÿ������L�/IM,��-9��1�#���X��%�d��0��5o� ���A��W�XrĜ����߯�_Gxÿ.�h�~U|�7݁�(W���X*c�͜3��� �ǅ5��ୋ����k�x�1Z��y�vы���y�ˇ �� ϊ���ߧ��t�6z�q�V�>�M�������$&�O��]9cꭗ,:���b�H)>�:%J��a��"�p��$O��yr���6SN[�8�����Pyw"�P�J��ARf�B?L���X��-�� �~Q���͢��nv��mBqQ��<3Z�Y�;ɢ
��/��A���� ;8P��&�x�,���9�S,��%.{gCB纹�x%V���S�`BVST�`�� ��[��w��r�>��z��n�Eu���d��)�ib�5Ȣ�a.�=�����,@Z�}��q�m'�Cxq(Bq�ZZ�,��k����m����D��N��<�6�]t,nF��rf�c*&c�@��fG��5��{m��~� �K��#���
W�韯]�Z2w�S���?��-:�&���-,���8����'�}*��:SH�r�L)�p����P$΃��n1���[��a���&N��N�:X��Ʋ1�'�X5�<uA[�QR��X?A�M��H�œΗ��q�fO��`��7��ޜ�۰U����[&Ұ����ė� �j�M������l<,� COq�+�.��܁A`v�!g��!���:�.�bj�NL~gh���WiR��p�(�5�6�%�XO�j�Fǆ,R���x��Ge8lC5u������x�XhО�j�2/P_�ᯟE��&�`tn��D:i{�,�Q�s!���6/+D��r��u�^j�]��'�U�#�k����}�H�v��bP����Hg���(�j��������]44h�mo&v���P��-{w*3�0����2�#%������ ��[�ߺ���Ʊ�ܴ2�H4G?�Ϥ����1J[��M	d��]Iի�cSK+�#q�F����,�j�U���:���K���Q��+��
{�����d
���
�&p�Ð�o� ƝIs ��1z���'ݰ�yO*�_��!�J�)<�q�[v���?&��_���ڵaiH����%JVv��}ǂ]����-� ����z��H`%�-p��y��ӫÈ��\�9\Bh����Brv�+�����r�H�4��a����۠f춲}�g-�r��=j�i?4H�;��I��&��}�`��x�Q���w�ů�Op�o
��x�!M��a��ϟ"z2t�bP�j�񝫇�Ǵ�ãU���������X�����nrOK�[���V�d�K@Ol�B�P���Z.�b�'�%]�qH�n��f��Tp:���"
���)ͫ3���2w�	��z-�)�$ m*��n�t�o
=ɼ�2�D�8�	��fܙ+X ]�m�(M�o��Df��|Ss�kg._t y�5� C�ŋ�M׳�+�i��7#^~oH��/V�����}_hk3�i�>����y��J���U<u"^&����>W��W������u4�Q{��Z�XM6|�)l��8��G�:�0� ���oTʕb��՜�a/
+��Sg�{%��]Sp�wQ�j͈�~!eJ�(n�4��4��ý�����2X�t(����d��@��ɤ��O��|i�MG�86��rt�+��
�j��_Ę|�&d�`���1$�ׂ�l�G�ꎍ�:N{Gt��P	3O1���Q.�1<]���SJ�����U=��R�N�͉�\Fϊ�R��w�o~��'���Q?�����y�ED��^���FV|�C,6;WT�D9�
 D	p���2�k9�����Q��)�0(�n'|�i�(kB�F�	ô���η�I�����x謬%hCA��8�	��/�v�
��6d�-�?�y��Ĳ�g��u��}����m�0�Ó[$5�ż4f���؇4Gg��P��!��3E��b2�=VDa�,ظ�^��Į "� �
�q�H��'�wk�?�B^[:
�����w0�k�uy4�K�{&�a�熩�����7�����r��L=��O����)Yr:�}�H?�=��Cd�je��4��Fw~c���59~��?Ie��I	����!s#�Ƙ���_��L�{w7$�k�6bcB�\��NF.+��tsR̥+3�
a�n3�BT"�K(��KD_R�KbX.s���?�_������z�ޯ�/���$���l`����b�����T���*�)��$�ֶR��+?C�u�G]<>?w�W��u.F~�hє�[�l~����F�����K_w$�\�g��D��aB%6=�
҂����PF�#Q�O2{.����$�ܔ�q�+�y,�!=2�zY�-R�'a򽨸���]	���tl�aЮ�$�1�toad�������^^��vNDa���C�)K9�ٓ�U#s�y_�ٸO�;�R���f����EAMﱘC
�(����xkQ�O��<)��S��2k�g.[�v��.]/��_��V-�Y�>��@:�2���d��,�x���m\��
E������cMO�Y~ڞi ��W��)8���4��Z|/�Z�f��f�-�A+v�]�$��m'J�gq�=)����5�9�P6j{K�P�Q5r�q�q�,��z�В:(������±Ŏ����(T_���Jc4�,h��;�yW0!�@���<tK6�[{�pЩt��?"�r����?2�l��ܯ���:�k��/0rs���D���br,"X��+��j9߹�7���J�{fY{w��fȗ�e߁�z��<z�4�q)�D�t�I"fdL�)�ݍ�ϥ�,�}�⑑���t,F ���u����1r!<:�Yg�R��JԵ>�����6�69K�)����ԙ �����zX��]Nַ�������)K�J�ټ[,J� ����;�}��Mw���W<���"밊)����){�F�9
�����wz�=�Ĳ�ŷ�k���Q���ͺ$S�و�6y��Ww|p�/[�l���W�&�|wK���[����T)�H��(��:��|U6=2���*�#N���[�_(���f�R����'�G�m���}�Z�Q#�nf�0��lV�lK�A0F��)�O�.���}f�.�ȧ#���H)B�$��da�h��� �&i��2+4�pE�N�����`�f��d���$��[̬ϹZǟ�G���DDs%h�ޚ���T`��2op\�5�]�g䕈	 ����rݖ��牢�W���ND�TRz����\r�r�R8���&�-z� �J�G��x�	��>@{i{���Xn�F���
��~��%�%��(�_8�d&���+��>�H��l|�js.Q�ȷ0�e賙�Iem(2нU�X�q~!���d=�-O����]M��g�9Y '^c]i�*�X�qJ�3��R��B]��o"�K��-P�ܒ��`���a��Է*D�;��u���M�m[�dZ΅��F����5k����sch�@C��z�.�� ���Oi��ۖ؅4.e�$&�B%������y�����u��R���	\�T^�j�a^�Qc��.��A�mx����4��ht}�hg�V��dGA�eK}Pk)Qu/$��R^?�2��q�D`tc���<�-��k���w&%�P����#��Yx���C�衸'��@�EЯh=�b>�g�/_�2���`�H���k��Prx[?m�&ѣ�eN5~��ˆ<�P�0<}��>��&��p���J��������p?��ݶ�ػV'dH㨛�ꕄB>���8T?����7o7J�U:.��	\�0�;
�V4Q{�jNRH����f�Ċ�0vJ�x6�Z�.���3ＡCYE�;P����ӛ���f�t���0 v-�����3��5����T�N�L�l\=K��ė�!<}�]Ne/ýý��o���T;��%�Δˀ2��R��`��L@;Cܫ��Pw���?�Ǐ��F�-"�k�B
^F�
.���v;V7�^��O��G)~i��.�M˾X���ݯz���v��A�Ψq��w/�w��l�㺍�_؜h�� ��P�V�f����yul��[t�,��y�IM��k��m�7b�o�� =��̓n�U}=�Z=��vӯ3|�F���$H�l��.���^��n RM6�Ʋ��ـ� 0�`<�؂n�ф���&�M�2h�@F�xsI�����;d�F־dGzO�>G/� ����|�z�d��ұ���s" ��t�L��})�n�a[)� ݡ� ��;2g��?�l���|"���z ~{�E�_��2�R�$�nS� �=�A�f8�`*���ܙf�I�(��s���h>��ok�[����]cj'����c�{V{��p��PK   �n'Y�T��[  �  /   images/ff38abd7-836d-491b-898f-03e44c25d606.png�P��/:JEE$GQrΈ 
C�s��� �Dp��38��Ȑ�D�"�$�����}�u�ޫ{_�{u���f�Z_�}qu���m]��L'!��5}��O�$Fz���'<n�xC �	��<yq�T��Quwu�w�x��ɩ�h�Z��ݾ�#'*)�,'!!#".#")+*+!#+".)#)�#'&!"!*!*�?k��M9݁�@un�ٺ�
Y۹���z@?
r�����5{�����\�"8C�&�)�d?�Q�s��WS?�
���w���CNX���_�_\���QXTVVVXDLXLL�!���c ���P�wRj�޶^N>N�n�߭m�}}����E�cg�_/�������=oaQ!����V�����������c�ŉ�A����Q�/@������ŇO����ދ����� ���0q�,�Oz��W�(��P/'��0p��G|	� �
[�P�7���T��������@�����a�ȧo����ek�?T���S���P�ǭ�Xs=�G�NI��Z�VF�F��A�^P�ABBPF�AV�Z\RRTJL\�ZJ�/Z�%�AI����\�pYI��ր7�c�w_ۻ�������?���f�w���GX�7��_�`e0R	�n ��7�z\��箻���]/'o'k7@���.�)�g��=�����D�p����j��g� ������n�c���u�_L�/�j	y���r' kiP�"B݈y�<�r��))�=lB�A�])��������{Q	�sx�4x��[8{��Y�K�LĻ�64��r�E$��WA����G��N��"1������C�� �#s
�_p����� Cy��oOҶV����)��A�!M������t������N}e���g̻���'T֜�05!^/1T�K�ߋW���Ӂ۱����l�'}-��*+s���j���B�Z��si�	uQ�0��G�`H��Nk|*����.�L_F#M7�2�]�vօ��-f��CEfu�A��s;���$�H���L�#�uA�]~Q��s���Ǥ���m�wF����}�sY�W�¹����K�dLFM���[�뱘>/o�Z��W�=,���R%�hf�r�F&��򥪳P5��U��$ۍ�9�N�X/��L#���Af�X˴U���s cA�c�GZz��]D#v�~��v��[_�W���}�z����0�\#�fԘŒ�E�a���]p����^�7�M�h��i�Ѿд��=0���7��)k�y�=R�W�m�1?�~�^֬.Q�`�s+X�"D�5���nqk9T}sȚ�s��PEEѹ��FH��ffgl���/��~p���Ɇ�C�v�ZBYH!������g�8��~��q�P�uX@u�OW��/%�L��U�Ʃ;��}%�e�nu&v���X�A�#��H��y�oxl�]���e��6N4,��:o�i|&z�(.��A�^s�x��Oz6K��`�|��3���/�_�$3mtY��wWR2�It��8�6d4��N�`�7�ߞ����	Vg�B�1Nq�M���d*�cY\/=�7@�u4�5�����싏���uݱ���z��0!�G i��^��6
�,�ی(@�c�:Xp�1��x3j���_�FC&���O�ŝG��-#M���t.���w��w�	��p�N��L3�1�(�»��_��{r8�92���8�p.�5���>�a
ơ!];?NA��C��D��YƇ�"���&0nG69��4e�-�Y����ڑ�ME�G���/;��PJ��#���Pw��pE�D��������v�
��wդ����E�c�C{�Z�n�g��t�N���ʪ]�S�n�`�@[q�fL�&Ŏ�NH�j�/���DC0ET�`&�.���]`%	�~�p�l�~ �u�N�:����03_��p�*��z$��Yv�^���K-���c��+�z09@[�c�?M�C �� ���!K=-�j<@b���d$���j�buʴ�%��ʧU��kd���� �oAdY��`t�4d��N@��� �Dt�H:�T!j��&rN�=]!�`� ,�=Z&,�ZOX&��2H��)P�٭*@�Fj��;���R"��,k ��t�O� i�S]N�)�r/�?%��O�X��A����K�oA��7��9��2��n/����?!s��P,�q$��9��*bJ���L���/�Ę\Q�P;A�s���g���9cJ0��I2�hQ��$�$Q9��n�!n2�%>g� 0[���z>�ݶJA�F���ez����O���SNL�*T*���i����?%����s�I�љ2���b�"�Na�:a��P0&G ;%�`���[��B4G��sTܔ̾��j�����b�}��������!~rL���A�
ު �P���k����A�y�L�L��0V���$>�"����-�:FL�����Z��I��o4��m���1�r�/̓�i׆�_���b�=��?'��k��� s����;����,z���;�I�{�N�_YI�h�Αr���ʷω�7<U�C	q1�[�(z���a�A:簪�p9���fM#�̧�,�y��t�Go��_��:�g�0���݌�}�e�FS>��۔�]��7�n%e^�&��np��������_��T����|�k}�@��b��$��ę,�A����e*�9���~�I���V@'%�(7s����x��{2}�M'���d�
nf����/m�����N hUj���k��D)��+�����*�$ tQ�ӹ�u~�r�?��ˏu+��P�V�ޘZ����|�b �Z% �y)��;�I�_ǎ<Ȯ��a�븄�K)v��ӑXdtS�?Vq�����{��������7SBx�7n�,s4�ƇG�iUɶ�'� 6�T�EΈe8�㕓C�N��hH�O�&$�B�&V������ a"��L��@)�|kP�*��v,L��>�u�hq%/K�g2�rL0��2�VZ�Qh���Eɪ�e�[���N�򾢑V`XRt���8��ۃ�_-&��<ٓl��w�-R$K��P9�6�K�}5)��(�.�����P����f�hfg�@��Y��,(�.��>�uYH"Y~D�e�h�x�����a��ߎ�Ǜ�0�Z��|;&#�~�"Խ[o9Ky�Y?�=u�#rǊi�*/E<=bh[&���=vn��Q�:k:4ұ65(����Y�����U�a�N)ב�m� a�L���eoltc�)|x��VՓ�������y7���Y~��2��7[9>�WJ�.�f;R�ݹ�f?`�Z�b��~zӾ���鏥M�q����ժ�~�iB�dL��+S2�Y��楬k��RF\[��{'���`NB̤%H;G��o�+L����WE?�ix��க虹�Qic�J�S���Ej�=dO5�|�DP���_����	�f�����.~����p7��O����χ �=�ƃ�� *���wI�1~���<u/w�s]�n���@{(��k�]��4�)�"aBi��Ԭc�qp��(I+�1�>���""LȾ��~ϕR�+7}|)���$_����-��@x�X���U_�ĮJry+()n����@]ݶ��qE�>1�ݐ��ۏP����y0��͟u�`⎲�	qA�\��t�KW�c96��l21���~ES�t�'ve�!J@~���B��۹ѿUl��RE��[��9̽�&
�\�F!�������.Z]5�n�XF��Gc/jdL�R��!t|Χ��˪"��R>�� �r,��E ΰ�"�*��`�����a�����جZ8%s��OK�Mm�#<�h���en��t`��,�>RH{_����ܖo��g��Y�%����\.�#��$�is��ލ�M2T��u�����y��6��8<nP������5ܷ�@80}[�FHC_rlBbB�A���8 �m3-��?d�y�4=� �syjA�|-�Wh_kw�t�d>�"��ԏs&�]bQܻ�K>�v'ɴ�}Z`II`�_�;-��=s��2�v:d7W*�M���{P֖�/����5�ޏ_ �G���uT��5n�LCC��74�B��	@4�iRb5J��6O�y����m���9 V�u���C��#�[�*ĵp���'��"U�P�H�S��W A�*�W��h���,YHlg�=`�^��?׎T?���F/����$���%�EK��|��Nz�/�N����c��|�µ�����8��]i�����i�	C�§�dN������E��� F�e��J}s9~��[��
��D��R7Pw�&B��Z�o�#T���"�X��<!L��"�������h�1��'�n�{��
qBf�?;��rd��'��C�Iƶ/(�/Z�V�%����ު���c:�C��0�8G��5s��9z��ߕK)�;v�>���Q�#��Je�
��n�ٺ�-l�q5O�����	m~�Cy�=B*9[�Uδ�n'Uc�Br6���ִ���J-"�}��|��>��M�7U�h��@_��֖�z`�uaׄMU������>����1�<�O�h�)A��V�E�:=�NO\��"L[�E���9���qr-��dw6Vr���v�d3�Q6��3��v�����ಲ< %f�[HW_����T~4�X���*d��J���(#�^��5���\�x��6Q�1A�1q;�wgW��~�0E�J=ް[6-�a���e�����n�"9�f���mø<B�!,�w��5a�fKQo_~�͆�`%�'�{}s4��)̓2��2��~t�L�t�r��Ȓ���A���EX�o����da���o�~W�)�Fc\��(^����T�Uʑ�v��l�%��L
(^h�K�5G&�xCIW��M�$�#�Ԏ����?�(e�e� h�4�
��A�6���Q(��v+h� 4�*<��%�~����<0b�ؕ��hw5ҧ���V��ځb�W*Y�  ����m��8�@'��0vl����F)�%�0y×K���	�=���I��]�R�@�9Io�s�2a!غQh�L����=��^PҤsd��(x�)���y��i�^�2w��H�
����E�h��X0�CL��ǌ�q	-LO�H�R��X&.,�P��jBJ�k�O� d�e���X�Zl�r�{V0�-���fj�;��'����d��ʀ��m�b�y�z���1Ec�X̓��l���$�#��H��Td�����k'�`u�T��X���sSDT/-�!�Ht�Փ�T��H7#���_M�[�+<�[�I'�k��������w�����w����`+�4r~'4Ē�[�iˇ]}�n�wW�����=la�y����؈h-;4�l��c\�°{�-��2��2x���H���&�wx7�M�Q��nr����&~>h%D����1����0�5�����ռqC�F{YT��^)a�	��Y���%��(���К��!T�@3r��O��Q���D��/m�.�/P3FX~"����gwM��;�d��-��� я�4�U,w�щ>o�J��=���<]�) �0y�&Ilĺ�1).�
 ĭn��^2��9+�X�r�?8�N�6|���?�73dl[s|�yş[�a�ɝ�gNҞ|��g�9��IG��r-O�T�(塪���+̍�X4�K�4�v3��^8�� B-J��G��{�}����Ghd��<����%��R�@6e+=��,�h ���h҃%��zܥT����GO�u?�ǡ"��jL@�\��{��/Q�]7>^�!d�jR=O�]�2�'��#%3���0{еD��8,�eg���*]�-�DI>O��h��ez��ж�d���g��(�i�6���;Tw�F�y��2֚f��h���q�W���W�R��%��xk�7)?8uKA�3�˒�X]`�<��>�ia4>'�sF�\�OB�)]��4�_�cVkU��|��#抅�,4u C�������bq�D(��tBP#��6R֌6�Q����4s�',$��V�Z�������� �p�(��z�S����Q�م��$�V�j�E������ B��Q$�1!�������PC����O<�i9' ���wy8��m��]@��q@�k���h©ԫ�����O���u���㤆�8�L�ȴ�M��45�H�� ��\�W���A&}x�������D��w������d�H@G@�0Y//ő~M�/�~X��_��#���5"�޽���]��.��!���14t���'�"��I�cc��y�`zV�'] ��vqP������˾�4�m��g��>+G�Ts�,��`���8c�R�1����CO`pꮫ�B��,��T��5�Ɇ>�9�4�-'?�]�<��%�S0z[\�#�u?�N(�f�$�L���B#��<�~}��D܏|�uq���50� ����ͩ[FtL�/��bb�˸��&��3@Sw��?i(��'3�����"���X�hT9�>y�ER�n�������m�'�Sq�0�jt>�
���|�P#[�kh�~�G0�1�������>�6�ꡚh���$	�`��p��yz�RUS8�ΒsRǏ�f��^;�9mȏ�b3)=�5�z+��4f{QA�`���{&�~�����AYP��H���m�{_�D9��A��X�h�M�/V/!�P$�+h�d�}{	���-چf� |��Pj&4H���U0�$OV�RB��_�T�ň���A�>$9n�Ȇ�yW�ނ������$x�I��a�қ-ֺ�%�ƆP�[�ǥ
���`���m.yP���Y�c?����D/�b�D��� �Q �i��c��(s!�`�6��a�r�*��CN�!T眪�i�J��/^�����@�n�T��[�X"l:�S��gx���issK���'�t�5�ф�W9궾�9�A�;��� �~S��c���� 7�ˡj�]`p��F��V6: �ݶ�$d�@��`���GS�����B��%��Q-���OTE�E��j��r����[7��͟�� +i{��	����keZ���n��R|��kKƑ����:ۅ/b�C�����Z�h�:r$� �ȱrN�$���w��	"j H����N�TX��ʐ��Ym-�L-�ܾ��Uq�� �4�`��`����L�XJs��B��<Zđb
�Ӓqx�=I�`|�e�3_<?{���7{fC������R���e]bI��jEjS��x\:h�|,�a�6��.ٙ��f+jS�Ͳm�۰:�g�=��B�x�땏z��y��+�wp�s4}���u��oR]���ʆ�_;���~���j2��q�B��x�3�t���&�P��`�/д�0P�hz/�-�5�-�O�iE��7�=0خ���g�1s7G)Mۋ�b~*��)�`! |Ch��I��hr���-1��N�t��"a�ݭ}�Mu�b��b����]�3-�!9�f�8�^��6�T���U�S�g	s����?�eN�#���	�W��
&������i��3(���ؘĪEª��g��
? �S���y�cȍU0����h�10*.���h\��'A�c@�v�m1 ��C[u.b���X���E�O��=3k(��r��Q�x9���@c'kb��[�D�x��3&�@|^��=V��ː�X�������Dt�	�U�9W�ꈸ^��H�: �Oz�I���`U9iC�m�-Md0�b"��#�=��dƣ��A��$�����|���1�B���+�T{�mͥv�6	�*$$ձ85�oerNd|M��(w+T�뛋�ʱ����	5��)[vM��`5����Z[��>,����k����
��A�� b]�?�z�K�j�e]�(f�� �#<�)�o��혾���h�J�l�c�1���6��us�MM��iT��1q;�é�����w�삪�zyz���]t*�>�C#�U{95��������1�o���r��l���� 6���R񯃽L6]d�N��͘�.������c=�ȼX��P. Ȁ<8l�:�	�Ѣ���;��n�}{Qbwv�D��5BCE��"�w��[�aɀI ߢb�z�8���O��F��=,��5�#��ׇ˷�^�/c�æ��=_TЯI��=VVn	�k�߳��S�����y\��zo9���C�3{���h�d�$4*L,S�mCr
JaK�y)��2
3yq�qk��'�2������K�E�W`rQ7��
ld�m�q�[�yK�^�����
���qz�3t�����M����u�·[u�|�e�b���C����O�0 �ӢХ���Gn�Z��E�\��N�h+�Ajw�ɊBʃxL�`Kߤ�rȿؤ�ϻ��&��wմ��|~�r�hm�,�Jֻ���&��#��&�)��5�f�ܗ��!� �~���!����/��G���U��樊_W|�֐�9���+}�g,��ԹwZzΏU�eee�ə�TχN9�C��C�I`�3�lٰ*��o˫킗�ƾyIP�/���V�'��`��C�o��ݻ�;ic��P�L��Ju��&e$?��o���?��&����)�H���]Fz�:�-ُ�}�
i����=��7�Ce��v��qW>�'_�#8 ����r~~����7��x3�UF�5�4d���y���5��=P���&e27:zLO}�\�X��ϔ���	�9�m2d�n�];�*���7h��;c�ރ�٫.H�p_�P���}�Sr��ʹ�
m�y/������B�����{��p���^��*�_���9V7i�ಜJ�zMu����%���+�4��SS�gMH5�.�^>L�d�y�z��t��+JԄ�x�B���V:+�l]7-�v�N#ͅf��KS�w��:�ͅ侞!�v�����\ oH�E\�.q��H�*3is�P��^�/���+�stu�"�
'>?Ӥ{����;��h�����耓x��k��t��^���Z��h���Z��E��@S�>l X���'�+:2��)6��Ahp�>�f���'��/�Pk���=A`ٝx�e��*c��֣,���&#�v3�$XtzMr�U�N-����ŕ�E�<�]Vcpn�`���"�i�Y�2�J�n�k�U)��tA�aJa�Y"<�W.�E��u+n(Q�����0G��������D�1VRk5_e�x5�]����X��Y`��3m;F�:B�ؕ�e�$�!�*|��/�@�q� ���X��K��
n���wz�x��g��?��Ix� �ö*��E�2~��<��Z�O�.���=��Voo��8ב� �*�]|l�^Akt�y�(����g��0�۝y���?�A�P���%t���8�m(�~=���*O��M��R�\�� ��uH����s��e.�UH`���������1�N�UJ�a��R�c$��64�}G������G=�wZ���8e��l!+=�����'�"���&��ȋO��y�3!b/�L�M��3�ǵ�ǌKp���vA��j��ꠕ�4�ܻ�5� �FB̑~����
�X6���Mrp���giER�����Uy�L(��/�"��|{;4�5=�l�\�l�����:D�W,-�X�t�r@#]w�&\�DZ-�Wm�����L��E��Ek��yW���Y{��{�e�B ���ŕ��LsA#�߹��p*�������TV�g,�Gҳ�x� U���6�ub��i�'�h%u���+�<�Zù	/��^Ű_pG�ɜ�a�/T�� M�<��]m�fa�baf�/�S�5�D�y��Jz<}�F�&\'=B���]��Q�~߯����#�3�"$�0��~���w�4V����ڟ� 8_
�FR�hʧ��W��Pػ��eE�Z$�d|-�s�����s�����m��t����ʏ�*�b@vR��{@��7G�	�Ey��L��23���1�+@��nD��V���L�)���t�@�����p04�3���Q��W6	w�[�$ٟ�T�B��xI�}�^M}XO8
qQ��@�:8H����{'(nKfw�l�K�,a7���8�ɋ��W�5I%�k�	�&E���=�ʆ�=Y��sT�Y�?�Z{D�1]�ֺ���6]WhS���]�7I��� �JL[����uo���^8151�m�E)cБ�h�����Y&A4~J���,[EZ�C�w���4��u�͂R��6;��Wah2��~��
`T�n�_i&���5>%F}=�߉�����`�� �oL{߾�s|P64�N醝������X{�Z3���u����WE�2�ݞr�ډ)��b&�������F�\T��AO>x5�`����ze��}�U�ʰT�(��U��w{e��;���	-�ޏ��7=���j�����~���
:=��!�?��X�V;��ȿ9n��DX$eH���Y�Q	zCà�I G�6�4������/���#l��j�A��μ|��Gk'��th�{{FΕ���9�j��/��;Wx��?_�6;~���-a������o[�7�85��OS�kn�}��n�����
8�z���X�P3��w�j���O.7�y�P�G����yj�|�i��0��t�.��O��a�Kk3/Dq�<q:���
�J#i���q��鬖p�s�������4BѤ_��(60G;��@3���~���/�;�6�/�������#9���W�;M�>(2ѻu���*�ȩ_���Qidhxg�g���.W�N���1�	�1L)뛒�7����l��m��z�R���B�d�Kw)30qz�m�w:�����5��V�1�PM���67���D,��_�+�~׻�|����d���#J �<�aa���_Ă,�|�ɤ�02�%���永�cy�?4BR��I�ܰ}cE�*F��<%��Ja�=�p���!�	l��KӉ��v�u
`h��u*-cNV��vP��I���a�IK�y��Q�.�D�cR'�j-�����b��i�4(�2�ǐ���jj{t���5%�p�G���
��GbR:>5�n<�Rą�߼��Gݽ�Oi��Nl�>�,�'�	ƛ�1x�9����_ߞ�i��	O��>�4�RS����Ó�&���ڜ���!Ws�����G]a��L�(A��;�4�u)�f�uiO���i6t$t��7�=��c�����WK�8����v̜~��w��0�=�!  ����_��}s��b��3��x��RE% : �=Q��1�`��T�W�Z3~�,�8� x��Ip[��Zp��P��hX��]��K9E*aKK�m+\�7_���}J�w���Gæ�<!�	�[M �vu"%�A��q��+��C�YHo���}���������0��\ހa�\I�'̵΢�����f�����q<�n��Y�s��k_���V{Wd*�Q˻9n�>���ס���jD����YD��:�[0��}��������bK\�if��yD 5�WS�2m�{3�@�}s������o����3`!"O�g��(�e�An<�/��~@�#���1�h����d���k��*m���o�o
�#�浅vH����q�ୂ�[�8�����:{�/#%��#nc�&��$�i�i.��S�N�-���5�s&�q֝�����s��}b����ʀ�`�r�%0���#��>��|�M9��[^0�p\�$:b�GK��J�|��i\�ҿ�>�Ku��j{L[���c1Q�.�@�i���D�\�
�3��1�_�F�$Y���I�v��?�_�m�F�à�n6^���w.�i�V�������XDVnNώ��d�x���ǳ�چYpˇ]�M�m�z>�ɋ��:�gE~`��N�.߰8��.,l��~�C��l���PBd�4��[��ȶ�_`K"�Wi�������K���\��S�a�Q��-ԁVn2�O����JyV��������ɀ�G�[Z�`�<5��-�m]i�eE��;���Ɲ�s��Ɏ����8�8?��1�P;%[���m����i��Ɔ��H��tg`6	��@��M��Ξ
��B���2eK���<�|?!JD��iT��p�@�޹[wg1�KZT�[+�cT��s12�����b�6�'�$6޽Ĩ�63��-�yo�|���d�弉��}�-7��re�vBě�;9�?�	w����,���k��������2��۰�u=����r�J��.��>
��LH5��R^|��)���������p���ŕ{�Cd���'�YG��o�@�h��ȹ��=��?��F���)'��R~��~�����I�%F%��iv_i$u�~�CIq0���HIj-yi�c��3��7�-P�gƗ>�R2����߽Id�/��Jz��֏��4&-t�I��j�S�Hv���X�'a<(A�#a�{2�z��ئ}�G	���0���H��5�f�����<��<����	H{�TY�Ͻ�3+O0�2D���D���hN �޾z�>�s�����o��{�4��uD?"�7`����ꣳ�7�:�7j>:��>b�O�(Pv���.�q,�= 4���ؐ;O�fy2�_���]5������;�5�K��g_ɋn�|���_��[��F�?Q1"5�>��"�%f�����Y�U[$ߵ�ΰ'�/�	0��ar�G����zA��@
�e��~��f_xg^G!BM)f�{�gf�yt�=\�iϻe�/��t�!Gx|����<4��4���#�Bt��%g��/�!M	����]���L��G��Z;��Ag��Q��c�I**z��-rb�&0K����~�4�n,2�z��Y�k2Xˏ����V�!s;t�h�F�y�cd��鮟$^��,��Z ���?�I#� �g9~ez�H��m&2R����ωn�K)�8hp����' �x�$������ʍ%3��[A�}G�����l�Q�r�ڠ?~�i��'Jj@|6�`�'�pK�a[���4i���5:�Uq�T����lS�`�lVǭ�E�<� �T����>w�ً6���dT����7- 5A�Ku1#���f���u���8�W-w7��Ay|�͏��O��6���8s����,��t<�L��(9�Zܨ���&)����|�M��4�r>��m?�ρ���7Q��z/�.Es�,+���%:��Qe��ڨ�c-���Qq���P��O� ?�&�α�ER[jӼif���W�H�"'0R�S�L�s�p�9*�9ʻ����P�3��k�2�Q%W�Ax��
�jg�M��:�.���?K�싇�~@C�^!J[
1����ߩ�J��@�./+�b�կj���*/�$��"h�k���������I
>~��|�M�kx����=g?%m�Zǝ��e���^g��A3���Z�������<oV���l		��ݏ���2�迊�]}FXTo��Je������{۞�y?�,�3C���+��42�/�}�y����Qm&�{"�ؙ�+��,n�9=�u����0�J��)�����_5TC��H�$��΀G ���m����5�^63!���*�h3,�-V; %+���u��r�[�pEQ��,1v&«k�pky��[}�?EJ�l�k�ݠ���:^z"��ῌCw�g��ui��Y��~��2%���G։v�F#ھ�x9UI��P�Ru?"t> �w\����L.��:��s/�����*��)Q�Nk��b^.x�I ��}}�-0f7�.����:j� _����.kw�v�)�D������^i��j��2�>�I�RW���\�s�|O¿�9Q����6�[�A���ф�ä����,'�L�����W9�u(��'��^e�j(.�U�~���l�`Pm}^��	Y�;���壻���p��ю1���r��`˩fk�E�<¨�a�VQ����߯j,�}�#t���,�04&��#9�>���Fa��Cѷ+�_(`�ӿRD3u�~y���)�\�c�p���+��G�R`p{ƨ��H���l�� ���#>[`y��V<�ʳ�>��3�����k��;η�pA��bߘ@��'_.iw����$���"A�hQa�Ez�O它CM7aN�*4�4՞߽�|�B�\PYϾsCH@���dӒv�0��2����@����Y�
���-V�>�R}S�j�^)�c��Q�ևl��u|�4��Z�f�Yj��,]��%'�6��Aq���3~P�N��v|aeIj�\�GV>�6勯y�+ִ��*�KS��5�|���*:z�K�t���� 0���-��(j�h�=�0V*`�^Q��cl֞'Gb�dФ�����ݕ�ޝ���]�po�mdhm�/���J@�b��\�=gE\�������;0�ec�! D]Ɩ�"�z[���uQ��huW�x�gōPK1Og�5_n�#'z�����hJ��}�𫯹�7 ��T� �ю�߲�f���H�ߚ[Tv���X8\���׃r="F���@ȼQ\PSwn��@��B���vit𙇒IG�"I#���
���5O��!("�`�覈C5��c�O����|��0�M�n�3I��.�ƷfH����)��*Bv��n��CQ�	����/�k����ۻ3g\��o����)�U~���'Wn^�a�e�f)�숎��PI���<]iI���H���L�%M˓�yn�h�.��ֶ�R�y���'/˹���4?�������	l{(�s�Ad5��ۛ��mG�z���%�;���\�M�J`0��3fNCQm��N��<�S#�Z;�(>���t����Ƿd���+�-R?u|	��n'$����I��E���M�o�H訩)���V]Գ����J��qɿ�h1'��;��Ks7.�5�j,L?2ɘ�ڸ$���5^w�"M����;��d�^�����^�jҿq���W���m���T��D本A��m��nyN��ReC)�����I��Ѩ[gB���V�g�%{n8i/���@�}�#��'!��A(_�)���k�\\oJ[[��p~*�`|+]�}�e�|Ư�3��@2gG��� S�[?�x���y���X��Pbb�Yq{9�u�ʾ�]F~\�P�:�MIA!�E�l��8��삹m���ٻ�=E�~{�ԛ�Y�3I3IhO��m��ylQ��K=�-����D��a���a�e��6Ve�ݺ�Թ�Uo�������Wm�=���L�iP�N]�g��T]4<�6o���t��q`nsN]�������{:��E=���oHz��T������s�i�i��`� ��'�Ҕ%�S�UNQN��پ}� ��Ŷ�P]��;���!f��E���[ưo��$�I�{q1�G��i������J(��g���Wޫ�~n#*�0��m�1���㷷���2k�8��+�W=T�}�G1I�S�J��}.^�3�F3�CQ�վZ�F�6~[Xܟ��Q���[V� ��X�T�Rг=0S�-���Ǵ����w>r�C\T�g�8WJ�W�"���� ?�uw�D�h�T&���F�ys���'������/�6�2��G3�g��.�p���ZU��1�� /�@���_�V<���������[B[~�r�r��T�l"û,�D�qJ�����L)k�U	o�^p����OZ�]o�<��o���LI��C��PM^D���ӑr��K�O���.A޵ݹ?��RVi�����&ZT�w�ͦ3�%�����o�pCa�h�x[?j?7{������;���qM�.�E��^��"��@��g����Q�p3��4�mCo��_�3X"���Dq��a�D�Lx�o�5T���v��_��qն���丛��X�e���	!6���r	�4P뗻3���	������4y��\̖�m�q�UB^c*�\c�%�i8:W���Fcō�خ�qD�Q��i�o
�6�?G�lr�CK�T�%*�x��1v}A��eu<�	��׿.��UciWsa
�+h���X:����Xe���ǟ�G�lgͥ�,�_��J�ұ�Om��G�M
��}�Z��J����'?:�q�H�Ahp��Uی�%F��aa�,�L�Ǚ%��\������Ϥq������/�1p��ǀ�&x}�3&x<L��a)�g�^�T�#���w�����T8e���7�Ǆ��M���]�����1�
�<S�d猴��cj������Ҋ�bT}���i�c�.1�	1-�C���-�q&w�
���g�vH��t�d���HN[�z0��[a�!��y�	3�#�|��U��{���]�L�'�K&�r��\�B�E	%Z���ͦZ�r&,��O����˾l=\��/^�V��}/�7S�Xڷ�y!�D.Q"�l}Ď^��pF�
�!�G5O�?��KMThM	�1�C�\��Wq���I',�9�!�%1�UR#G|�x[�+�v?��#��(i�$������x��F���C>���6�[+�-���W����vo��������m��>��P~�L��"!��gz${n�+3��,�������S�tJ���z��z��\��|T�����nZ�WRc��*r�͂-:Jպ�|����d�ߞ��-d����	�,�릳&U�Ǟ�����E�g��,����7���k�z�C��j'"%+��~	_a@f�%���U�DT�Yw�@ɥ~?a�E]��j�P��FA8�sU�ml�
M0��4�tx0��ڍV�������g�3�E���^�t��ܕ�/rd�ޏ��Y�E����[߸���̀��X_�"�[��?k;f���N��8�"G�yf�èI6x&`�?�7s!c���
��$9qEՅ�:��-5fE�d��f��ӯ���C���g�����nMuza��{&cψ��D��B��x��	��}۫�{�R?�Z�/�
`�u �	q������BO��Xf<>�%�����sD��I& ��]���~���μ�r]�����w5!Kя$���b��7�Xc/���R�k?`�C^ ���=��t�o��h�c�5T������E��� ����}AXi"�_+�(�`�/դy'f�|;�^���b�мn�*9Yz+�%�j��=P*�/s�sRg��R��"��T���r��kq�if�����y���F�x{�W��r�w��� &�����chQ�+�ZX'Ë$x��X�&������[�.�xKDE��sp�y�A-_m���>�Y��ع�QAi��I�����lk/��P��zYzu=�3�����Qt|����:ūK;�8�s�~�v�i&\�/Y�s���^	g�4��{��K}�oLln����۳���CE}�6�s�!{�
��l
4�G(M�����⭹��������; O�9��x�޶zn�Z~�cc��?R	��S�g>�qÉ�I�����Ͼ���"Y�+<S�	���+�+y{o��n�<��3�̭���94Zd.�-
�9'K���_�B�G�	���n�~r˙�0݇4.�ٮ?2��^6吻,���Z�!��F��픟�s�تׁ�2�/�fcCS�!Gg��@��
��eܕ�s�Z�K���w�@���&a��c�u�?����?t�u�hn�P��`�T�t�.�<F�ъ�վ���G$��D���n�p�:Q���Gn�4��3�rjD��$�(�%_�[�c�v��?�͐3�@�+�Ȗ���3X�Un#��j��áܾ��)���D�A�H�&�T'�#M��b(1n���\�Lr�s
���Δ;9hj��Ȕ\r=H·�}��<��|�~|�����~�^k�u�k���z��3>o��Ͷ��=�؅����Y���5��VWп�=�Ϛ_�8A��G��''�k�4h��ޕ3�sɣ|Z�b'�3�z�Q�;��s(YLh'ϸ؈K���!�O6���|hB�u�,07�Iv�6Bg�7�,���&����f�I~
�ćn�^BSDc��{�B�P�@̐���^��D� NCKy��g��B������^@��	m��V�L�@w��"��E��(~hn�+���1��K1漢�^�s����Ca�;L�,�>�[M�*�ٜvԙ6��b��J��e��d<f�Z)�ɔo��_ُ�л}�_]9���H��WR�S����\s�����&6��ΰئ�}�q=��ɳʎ�S}�F��� ~G���(�\6����S��Ɂ��М\�Hǫef���bn�It�v��B�U��|�Q���PÜ{�X��8�F@��L&�k x��i�B
\�^^Q�Ԙ}~C�ŊhPm*�!MM*`��t�� �M�̿Y?��TeL��`�dsJ��з7����"�#ð�!ÊT��� ^7#W/�084�DQ�;E���tL� ��)02�1�چ����c��\G�� W�P�� Z�)�߹KB�kQ:�V��r�R��j*��ؿ`3$K�ړ"��)}�rEC@:Q?p�f�p�����	.��Q���@FH��s��͊�ƣr�p�;�g^���c��lQ	V�p�k�W Օ��$�,G�*6�.�P��ϔ���g)�p�k�)�L���w)�`Cq���-<ό��uH�j~Y_㗕�!�31�,r�����쫻�Υ,׭�^r'��E=G�ǒO�v�܄���&t��z.֜⭹}�M��mB���
դɵ���Bߑ����_X;%����y�"3��-��A
-PFt>϶��Z����d� , d��~%<pk�^���7�]�FS<�q��׻���K�I�2�[l��<��>R�[��WEE��b�^��߾����>�"~�(�<Y����|q�o�>:���{%�ǧ+�-,S�?���dj��?�Ȉ�$t_h�C:��z�^)0�}�gp���{Z�=p�{f^JGG��b�L/�P��~�Z�j���F%��«Eu�w9���_K�}'����oB�odp������ًwwבּ�s�a�}oԭ���2����q�C�Rf%H�����w�y�q���E�'| k�zP!��nw=�J]�%YԚ�T��`��r8u��	z�KU.�x	r�gaM�F��]]���:�w��2X�	)�JA��T���k;�(�*\�U����@�|S?��nCyw��;�xJ�{m���{�E6��r�W؆���wƑ�,�@�wZ�����5E�௾����cJ�d��zfjQ`RSU�f2�mG~��،� ��`r\0ս�\�@�O�;�'y�䷂�ތ7�9�-��lD˃M��t�P]cD�����.��=�$u0d���A�\� �L�w����^��T����*����3Oj_
#�v�C������~�.�gFޯL�ɱ��VF\7=�0 ��ᖬ��g̒�Ï�E��E�ܝ���yLsX,�td�Om&�%;���
,��.��cS���0����N���b'��h]7{A�@8JQ�ۉ�/Bȇq?�'�:'�(��3=�|H�)>�����,��{���_�MY��­׎2�����ڮ���E��NA|�BZy nG�}�%`���:�@�PZo�\�n���K~��̼`�U1������l�@3ĻDgT�����cI�p��kzc"u���V�x���H9����u���B��ⱞ��J�<w��G
^�w�S�����ZA��/&~�`-��V�J#wR�k+w�&���Ww��	 i�>�9��d�# zͮa��U��	��Jt;ݰ�'��lx%Z��{������9O0��)�"|�ʆ(^EOW���Ã�����[�!q/���k��`�������/ګ��|+�?]I�gi\�
��M),�`�}���@�5�Uw{#J�
�͈�'��tO@�d�/�c-<�!El|>��+���"%*|�< ���,��J[� ���޹6oK����x���i՝�l�=��\��'9�Y��#Z�!C�7Ӯ�(�vQ�o��U�ۧ&8ZtٚV��6�?#&O��%Q�)�~n�¢�� ����`�x��RI�o��&�I��ljo-FN�����ј؏z�Ѯ�c�/OhtS��J(��]�r	�0��	��ֈ*�8�5�u��Z
���3�sv��O	�u���/Sys�?�l�V� f��3�)<O��v��N�e�o��Ua�]��ּ֟MJ��@�`�Wa��]��!�h��餟c=t�F��5ؤ�:�l.6�2g�|1�:�e��:@���z��U"%n$��u�����s �l���zO��6.�T��N�,���8�p�+���C�n���,�pGi�"����ɇv�a��-�6҈"�f]l�]�Fk�������F���mf3�zR#���Eœ3�7/��m�-�sO���7�^�-9f���;{��n&�ωl���h�ݝ��	��A���*H��4��f�ohrjbA�:6F��ѡi�b$��L��ԍ���+>��GBLJ�Қ�8��moq��c�4.�㶳��!z��Z�wa@=��`|�AG��P�����Ora��؆ޅP��s. r�����/������H%X��%VOJh��~5��Ԍc%u%�$�No{)�����̷�i�C�|U����/;H�K��M��d޺��b(���{�e8Ï/LShͱ�|�>�6���?Ib9����U���e��ĵ��3�~D xS8��UL�bS����S^�H�,���%�\�*�����o�j�,�l�A��
��=h�Z�I��ƌW�N��i���V�c���Q'���u�=��W�@���Z�lt�פqL���
��۷�c��I�K�Y��$��RU�T)*�ʡ��9��ں� ���{���h����'�p.,���c^AW��/���[�� 3މ��-����8ө���zJ!$���j�D�"3���&����m����K�qLQ��f�����Õb9�0O��8�,����k��7y��	�?�.����g�+��pb�Ǧ��!ei>�^���j� M!9�N�~� WR��0ʙ}]XK��Q���f�HA&��[���L�% ŇX莇�Q$`Q g}A����I�.ͧ�Ưz�fSW�N�m=Ȱأ��,1�տH�\��p̎�zF�׍�p��2n�mCO��z�F������#	��IaU(�hI[]UIvX-�J�9���ݿZ�������e~���X����.9ѻ5���+�S0�EЇ�^�	�ӦPL EH��N���_���[I�J�,��r)��.�ᬕ���� f���QR�6�O�BH)O�J�-N�Z"g{��s%�M��\�zsGI*����=m6�����Z�| |���fz�De@�-�ܝ��]�S+�I�Qzs�[�^@���U_ҹ$��yn���ٜV�c/�}V��m���Y�z..�z�E���7����$�2!L�'s����J�~����_dVNG���Z鴓b��W�~�Yߞ�&��
ࡃ5�9)َ@η��jAH|}�`�̩~�v�.�:�ئ�8{���1R�,頍Z՚|W��١�����o<0ҿ�� }��S��T����m�A�K�w݋$���D�[J����؃�[���Ţ�d�7�>e�9OW����~4ueq��� ���}s���y}*�����Plo���"z5��g���O���{s#ʗ�6R��mĕ���ۗ����A]l��m;u,�lC�5�O}�l)DM���O��B���C�AL�k=ۙ�جC�v��M������2KT��! �@f��V�v*�Az�&��|C,�'q�:sg�� .�5Fޛ�A��0�gu���F�zv��c6�A���Ofp*=ǳ@���?88%��C�\�yv�����c�>�����S��㓞V'��^�W�kT�ۖ��wC�j�h�G)t�짔�B��G��SF��N�4����d΁���$�>�ʧ�w�/��Ai	f5�0&&�N���5��j;�g��^�*�0M�4L���p��ޞ��CةL�&�	�]#3\�8'�Y�a��l����sRg*����FX�wg�ޭ�-��KP��^	��槚i>��:��J�Q���#@t�c�4�jq��`+�-"��&HtG���?��}N��8v��\���j�v��z�������^��v�n2�h.dfYD@�GZ�,|�F<�t��Np/��32&�0}ó��#��a��3��,I���>�ؗ �L=f��:Р4��^����c������J^r����KK����rN89�c*��n��ߞO��@z��1��t� E�e�9%v�p�渪�X�=;BW�=��t��'��E��8�L�&=ڞ	)�B%��j��9��������b�wݧ��%!�b�	c���+�N��ANn�0<�:�h+A_��ٿh���$r��rB����E=�3lٖ����}nC)�m'��R���4Wnq��ot��9�Z8�d.{?\s���|�`x䝝w��dV�g����É��8�/�#3ZR9&��.��c�$C��I�0�A �R':�!*��]�T2228�_%I��$�������}�3厁s���JjG^j���:cc���h���+������m�i�>��0��B?C������=22R�3���g�`����:LcE�����WIW[Ơ�,�ءH#��,��4ϛҊ�M��zvZ�:��+AN>�����F����֠:�{���%c̊j-�S��m��˘?ׯ��yjm�b&zZ�9�=����Ĳ�:�$�G���o��/�履��PbHc/Tr��NCBH���p�C����y�h�=vn-b��I$�%
���r�r����a��_(eÚ���g�An�Ao��3����yƴ��Ę�(��J:,b9�a
y�.��6�Ixն�툝k�*�y@x��x�ɘ�a�5�TX�r�+����o+�型kFz�[����4mI����6������ƭĊLS��/���}]l��ab=~u;�n�]-Ñ��F�b6��Y:yd�UlJ�My���)mg��TFɌ�,��V��ڐ@���Xd���z�N�L���>��[����d����֚��e#�;�e�m�AqƏ>��fꨞK�Fs/��^~�!g���Rx�QԨ\�����+h�QYȘ���Y�r�������]�4��T�~�)6�5����xr1r�t̛EUF:�hZ/�zm?���yY��H��/�&�˼��2�[ɚ?�9��i����F��7�ڏ7��� ��f~|���%�/���M����!����@�凐�W�l���.��
����jv�z���PK   �n'Y���k  �     jsons/user_defined.json�Y]o�6�+��6�x�ͼIW[�"N�CQP�s$W�A�����iKK�����%��<�~0��헵��w�~*}�j_��[�n���4����.�n�G��?�8s7ݻgM���]����{Ô�����������ַ��Κ0������㢧<y`<ڶ;��Wx57E� M �K����K)��YŞ&t�7E[���l�
�-�����\"B�I��� �F�e��e��
߫��^�Aj� �,LĕL�O�|Yz�}|��]���؁���O�+�=>]W�i������ݜT���}9nV��s��4�S��켹��w��a�wu�y�_U���m�k��M7��T��j�w��ex���1�ͫ��nZ|�q�W.���Wt�u�"p>�k>
�j�����Qx��^�T����<B�:*Ǥ�/�(����0wƒ��(�����Ne2:�����+#�NF?E���MF���Ё�"Y��?G�m<K���!�+���<�r\�{z�Za����l?6-��U�&��|y1N�d����lAl]P�
���s��{��{�07F��+aT�MS'Q9�/�9M�;X����ǃ��*#��',�X���ڦ��{X���?�a{�t� 1��L&���v�P�+$���x�[ HT���0t�c�L&������KD�f� 61�~�O����.���J���b�`O*|L!�Ǔ2ݓ�{'k�N���/�/�F�j������f��mշ48�hn�M����c���~lu�_����ٹ�z}����}��O�lmf���T�#��N1b4+�ȱ�0�a�dV���i>��ќ�`�@�������g$�>/��k��KX���jo_�3�,��%��LYI��ʘ�}���L�Ƌ�8B*�1sc-��<�r�s9|S]�nu@w��B�P,4Q�"�B�
����8D�2lU�N��us��Z�}2�����a}���8{w@�b-VOڠ���j�3�U���2՟O�90���@
k�Њ8k�i�5�A鱩�t�[^��r��zt���{GK-��.a:Z�����ָ���'���F�$�����%���� �s��!�ь@�E���,�#��.��4@q2@A���t2������L��LͰ#�l���n9��X2�~��(����@53E�yF͵�rI��c�ݡ���zw�N�pgU9F{�:��5n&x����_Zg!pq���
9-��X�^�)q�"���k�1�)^2Lq芜It�*s�ȀK�u��8�����ð�p��Ufp�(4�4c����B�������Җk���Ǯ�-�j5{�T������7M�����aWGU�Üz1j-TnA(MArk�%+��VY�`�ﻓDVi9Ӂ��Q"�g�+	��]HW.����NPcA`�n�t�c�C*Lq�v�ӂ�<>�����w���\�q��<�`y��SV��̰B3�����*`� �b�.�~�*=i�T��*fj��2�dpA��	V��c�f�Gm��Y���֭v�=_�a)��>�}0�us��>�x�����e����v���w=y/���8]����~O�^����=�,�D�^�X %b�*䬐\��l�L����PK   �n'YQ��  �b            ��    cirkitFile.jsonPK   �n'Y��(��8  �8  /           ���  images/12674a71-c981-4176-a988-13f1272e71c5.pngPK   �n'Y8�w���  ��  /           ��!Q  images/54656ac2-7b78-4fd3-b315-813e86bdf352.pngPK   �n'Y�?HU!  B#  /           ��m$ images/585092fd-6de4-462f-8499-92296fb2c536.pngPK   �n'Y=��� Ѿ /           ��F images/732af9df-f9f3-48da-8e69-a852eebc5446.pngPK   �n'Y�7}b  ]  /           ��5J images/7f5f08f4-fdda-425c-ad26-fd4aedde5760.pngPK   �n'Y腸��� v� /           ���b images/a03bdc4a-b433-4a71-810a-a5f1c0469152.pngPK   �n'YXs�銙 � /           ��)	 images/cf59327f-2b20-4f20-97ad-1ec426c5b43a.pngPK   �n'Y��T�Y  I�  /           ����
 images/d8e70382-63d2-4b8d-b385-7bc04a585f98.pngPK   �n'Y���n� 6 /           ��� images/ebd5c09d-583c-48f4-aaf0-071f49184249.pngPK   �n'Y�T��[  �  /           ��* images/ff38abd7-836d-491b-898f-03e44c25d606.pngPK   �n'Y���k  �             ��� jsons/user_defined.jsonPK      $  ��   